// system_acl_iface_dma_0_dma.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module system_acl_iface_dma_0_dma (
		output wire         dma_irq_irq,                //        dma_irq.irq
		input  wire         dma_clk_clk,                //        dma_clk.clk
		input  wire         dma_reset_reset_n,          //      dma_reset.reset_n
		input  wire [31:0]  dma_csr_writedata,          //        dma_csr.writedata
		input  wire         dma_csr_write,              //               .write
		input  wire [3:0]   dma_csr_byteenable,         //               .byteenable
		output wire [31:0]  dma_csr_readdata,           //               .readdata
		input  wire         dma_csr_read,               //               .read
		input  wire [2:0]   dma_csr_address,            //               .address
		input  wire         dma_descriptor_write,       // dma_descriptor.write
		output wire         dma_descriptor_waitrequest, //               .waitrequest
		input  wire [255:0] dma_descriptor_writedata,   //               .writedata
		input  wire [31:0]  dma_descriptor_byteenable,  //               .byteenable
		input  wire         dma_read_waitrequest,       //       dma_read.waitrequest
		input  wire [511:0] dma_read_readdata,          //               .readdata
		input  wire         dma_read_readdatavalid,     //               .readdatavalid
		output wire [4:0]   dma_read_burstcount,        //               .burstcount
		output wire [511:0] dma_read_writedata,         //               .writedata
		output wire [33:0]  dma_read_address,           //               .address
		output wire         dma_read_write,             //               .write
		output wire         dma_read_read,              //               .read
		output wire [63:0]  dma_read_byteenable,        //               .byteenable
		output wire         dma_read_debugaccess,       //               .debugaccess
		input  wire         dma_write_waitrequest,      //      dma_write.waitrequest
		input  wire [511:0] dma_write_readdata,         //               .readdata
		input  wire         dma_write_readdatavalid,    //               .readdatavalid
		output wire [4:0]   dma_write_burstcount,       //               .burstcount
		output wire [511:0] dma_write_writedata,        //               .writedata
		output wire [33:0]  dma_write_address,          //               .address
		output wire         dma_write_write,            //               .write
		output wire         dma_write_read,             //               .read
		output wire [63:0]  dma_write_byteenable,       //               .byteenable
		output wire         dma_write_debugaccess       //               .debugaccess
	);

	wire          modular_sgdma_dispatcher_0_read_command_source_valid;    // modular_sgdma_dispatcher_0:src_read_master_valid -> dma_read_master:snk_command_valid
	wire  [255:0] modular_sgdma_dispatcher_0_read_command_source_data;     // modular_sgdma_dispatcher_0:src_read_master_data -> dma_read_master:snk_command_data
	wire          modular_sgdma_dispatcher_0_read_command_source_ready;    // dma_read_master:snk_command_ready -> modular_sgdma_dispatcher_0:src_read_master_ready
	wire          dma_read_master_response_source_valid;                   // dma_read_master:src_response_valid -> modular_sgdma_dispatcher_0:snk_read_master_valid
	wire  [255:0] dma_read_master_response_source_data;                    // dma_read_master:src_response_data -> modular_sgdma_dispatcher_0:snk_read_master_data
	wire          dma_read_master_response_source_ready;                   // modular_sgdma_dispatcher_0:snk_read_master_ready -> dma_read_master:src_response_ready
	wire          modular_sgdma_dispatcher_0_write_command_source_valid;   // modular_sgdma_dispatcher_0:src_write_master_valid -> dma_write_master:snk_command_valid
	wire  [255:0] modular_sgdma_dispatcher_0_write_command_source_data;    // modular_sgdma_dispatcher_0:src_write_master_data -> dma_write_master:snk_command_data
	wire          modular_sgdma_dispatcher_0_write_command_source_ready;   // dma_write_master:snk_command_ready -> modular_sgdma_dispatcher_0:src_write_master_ready
	wire          dma_write_master_response_source_valid;                  // dma_write_master:src_response_valid -> modular_sgdma_dispatcher_0:snk_write_master_valid
	wire  [255:0] dma_write_master_response_source_data;                   // dma_write_master:src_response_data -> modular_sgdma_dispatcher_0:snk_write_master_data
	wire          dma_write_master_response_source_ready;                  // modular_sgdma_dispatcher_0:snk_write_master_ready -> dma_write_master:src_response_ready
	wire          dma_read_master_data_source_valid;                       // dma_read_master:src_valid -> dma_write_master:snk_valid
	wire  [511:0] dma_read_master_data_source_data;                        // dma_read_master:src_data -> dma_write_master:snk_data
	wire          dma_read_master_data_source_ready;                       // dma_write_master:snk_ready -> dma_read_master:src_ready
	wire          dma_write_master_data_write_master_waitrequest;          // mm_interconnect_0:dma_write_master_Data_Write_Master_waitrequest -> dma_write_master:master_waitrequest
	wire   [33:0] dma_write_master_data_write_master_address;              // dma_write_master:master_address -> mm_interconnect_0:dma_write_master_Data_Write_Master_address
	wire   [63:0] dma_write_master_data_write_master_byteenable;           // dma_write_master:master_byteenable -> mm_interconnect_0:dma_write_master_Data_Write_Master_byteenable
	wire          dma_write_master_data_write_master_write;                // dma_write_master:master_write -> mm_interconnect_0:dma_write_master_Data_Write_Master_write
	wire  [511:0] dma_write_master_data_write_master_writedata;            // dma_write_master:master_writedata -> mm_interconnect_0:dma_write_master_Data_Write_Master_writedata
	wire    [4:0] dma_write_master_data_write_master_burstcount;           // dma_write_master:master_burstcount -> mm_interconnect_0:dma_write_master_Data_Write_Master_burstcount
	wire  [511:0] mm_interconnect_0_pipe_stage_dma_write_s0_readdata;      // pipe_stage_dma_write:s0_readdata -> mm_interconnect_0:pipe_stage_dma_write_s0_readdata
	wire          mm_interconnect_0_pipe_stage_dma_write_s0_waitrequest;   // pipe_stage_dma_write:s0_waitrequest -> mm_interconnect_0:pipe_stage_dma_write_s0_waitrequest
	wire          mm_interconnect_0_pipe_stage_dma_write_s0_debugaccess;   // mm_interconnect_0:pipe_stage_dma_write_s0_debugaccess -> pipe_stage_dma_write:s0_debugaccess
	wire   [33:0] mm_interconnect_0_pipe_stage_dma_write_s0_address;       // mm_interconnect_0:pipe_stage_dma_write_s0_address -> pipe_stage_dma_write:s0_address
	wire          mm_interconnect_0_pipe_stage_dma_write_s0_read;          // mm_interconnect_0:pipe_stage_dma_write_s0_read -> pipe_stage_dma_write:s0_read
	wire   [63:0] mm_interconnect_0_pipe_stage_dma_write_s0_byteenable;    // mm_interconnect_0:pipe_stage_dma_write_s0_byteenable -> pipe_stage_dma_write:s0_byteenable
	wire          mm_interconnect_0_pipe_stage_dma_write_s0_readdatavalid; // pipe_stage_dma_write:s0_readdatavalid -> mm_interconnect_0:pipe_stage_dma_write_s0_readdatavalid
	wire          mm_interconnect_0_pipe_stage_dma_write_s0_write;         // mm_interconnect_0:pipe_stage_dma_write_s0_write -> pipe_stage_dma_write:s0_write
	wire  [511:0] mm_interconnect_0_pipe_stage_dma_write_s0_writedata;     // mm_interconnect_0:pipe_stage_dma_write_s0_writedata -> pipe_stage_dma_write:s0_writedata
	wire    [4:0] mm_interconnect_0_pipe_stage_dma_write_s0_burstcount;    // mm_interconnect_0:pipe_stage_dma_write_s0_burstcount -> pipe_stage_dma_write:s0_burstcount
	wire  [511:0] dma_read_master_data_read_master_readdata;               // mm_interconnect_1:dma_read_master_Data_Read_Master_readdata -> dma_read_master:master_readdata
	wire          dma_read_master_data_read_master_waitrequest;            // mm_interconnect_1:dma_read_master_Data_Read_Master_waitrequest -> dma_read_master:master_waitrequest
	wire   [33:0] dma_read_master_data_read_master_address;                // dma_read_master:master_address -> mm_interconnect_1:dma_read_master_Data_Read_Master_address
	wire          dma_read_master_data_read_master_read;                   // dma_read_master:master_read -> mm_interconnect_1:dma_read_master_Data_Read_Master_read
	wire   [63:0] dma_read_master_data_read_master_byteenable;             // dma_read_master:master_byteenable -> mm_interconnect_1:dma_read_master_Data_Read_Master_byteenable
	wire          dma_read_master_data_read_master_readdatavalid;          // mm_interconnect_1:dma_read_master_Data_Read_Master_readdatavalid -> dma_read_master:master_readdatavalid
	wire    [4:0] dma_read_master_data_read_master_burstcount;             // dma_read_master:master_burstcount -> mm_interconnect_1:dma_read_master_Data_Read_Master_burstcount
	wire  [511:0] mm_interconnect_1_pipe_stage_dma_read_s0_readdata;       // pipe_stage_dma_read:s0_readdata -> mm_interconnect_1:pipe_stage_dma_read_s0_readdata
	wire          mm_interconnect_1_pipe_stage_dma_read_s0_waitrequest;    // pipe_stage_dma_read:s0_waitrequest -> mm_interconnect_1:pipe_stage_dma_read_s0_waitrequest
	wire          mm_interconnect_1_pipe_stage_dma_read_s0_debugaccess;    // mm_interconnect_1:pipe_stage_dma_read_s0_debugaccess -> pipe_stage_dma_read:s0_debugaccess
	wire   [33:0] mm_interconnect_1_pipe_stage_dma_read_s0_address;        // mm_interconnect_1:pipe_stage_dma_read_s0_address -> pipe_stage_dma_read:s0_address
	wire          mm_interconnect_1_pipe_stage_dma_read_s0_read;           // mm_interconnect_1:pipe_stage_dma_read_s0_read -> pipe_stage_dma_read:s0_read
	wire   [63:0] mm_interconnect_1_pipe_stage_dma_read_s0_byteenable;     // mm_interconnect_1:pipe_stage_dma_read_s0_byteenable -> pipe_stage_dma_read:s0_byteenable
	wire          mm_interconnect_1_pipe_stage_dma_read_s0_readdatavalid;  // pipe_stage_dma_read:s0_readdatavalid -> mm_interconnect_1:pipe_stage_dma_read_s0_readdatavalid
	wire          mm_interconnect_1_pipe_stage_dma_read_s0_write;          // mm_interconnect_1:pipe_stage_dma_read_s0_write -> pipe_stage_dma_read:s0_write
	wire  [511:0] mm_interconnect_1_pipe_stage_dma_read_s0_writedata;      // mm_interconnect_1:pipe_stage_dma_read_s0_writedata -> pipe_stage_dma_read:s0_writedata
	wire    [4:0] mm_interconnect_1_pipe_stage_dma_read_s0_burstcount;     // mm_interconnect_1:pipe_stage_dma_read_s0_burstcount -> pipe_stage_dma_read:s0_burstcount

	dispatcher #(
		.MODE                        (0),
		.RESPONSE_PORT               (2),
		.DESCRIPTOR_FIFO_DEPTH       (128),
		.ENHANCED_FEATURES           (1),
		.DESCRIPTOR_WIDTH            (256),
		.DESCRIPTOR_BYTEENABLE_WIDTH (32),
		.CSR_ADDRESS_WIDTH           (3)
	) modular_sgdma_dispatcher_0 (
		.clk                     (dma_clk_clk),                                           //                clock.clk
		.reset                   (~dma_reset_reset_n),                                    //          clock_reset.reset
		.csr_writedata           (dma_csr_writedata),                                     //                  CSR.writedata
		.csr_write               (dma_csr_write),                                         //                     .write
		.csr_byteenable          (dma_csr_byteenable),                                    //                     .byteenable
		.csr_readdata            (dma_csr_readdata),                                      //                     .readdata
		.csr_read                (dma_csr_read),                                          //                     .read
		.csr_address             (dma_csr_address),                                       //                     .address
		.descriptor_write        (dma_descriptor_write),                                  //     Descriptor_Slave.write
		.descriptor_waitrequest  (dma_descriptor_waitrequest),                            //                     .waitrequest
		.descriptor_writedata    (dma_descriptor_writedata),                              //                     .writedata
		.descriptor_byteenable   (dma_descriptor_byteenable),                             //                     .byteenable
		.src_write_master_data   (modular_sgdma_dispatcher_0_write_command_source_data),  // Write_Command_Source.data
		.src_write_master_valid  (modular_sgdma_dispatcher_0_write_command_source_valid), //                     .valid
		.src_write_master_ready  (modular_sgdma_dispatcher_0_write_command_source_ready), //                     .ready
		.snk_write_master_data   (dma_write_master_response_source_data),                 //  Write_Response_Sink.data
		.snk_write_master_valid  (dma_write_master_response_source_valid),                //                     .valid
		.snk_write_master_ready  (dma_write_master_response_source_ready),                //                     .ready
		.src_read_master_data    (modular_sgdma_dispatcher_0_read_command_source_data),   //  Read_Command_Source.data
		.src_read_master_valid   (modular_sgdma_dispatcher_0_read_command_source_valid),  //                     .valid
		.src_read_master_ready   (modular_sgdma_dispatcher_0_read_command_source_ready),  //                     .ready
		.snk_read_master_data    (dma_read_master_response_source_data),                  //   Read_Response_Sink.data
		.snk_read_master_valid   (dma_read_master_response_source_valid),                 //                     .valid
		.snk_read_master_ready   (dma_read_master_response_source_ready),                 //                     .ready
		.csr_irq                 (dma_irq_irq),                                           //              csr_irq.irq
		.src_response_data       (),                                                      //          (terminated)
		.src_response_valid      (),                                                      //          (terminated)
		.src_response_ready      (1'b0),                                                  //          (terminated)
		.mm_response_waitrequest (),                                                      //          (terminated)
		.mm_response_byteenable  (4'b0000),                                               //          (terminated)
		.mm_response_address     (1'b0),                                                  //          (terminated)
		.mm_response_readdata    (),                                                      //          (terminated)
		.mm_response_read        (1'b0)                                                   //          (terminated)
	);

	read_master #(
		.DATA_WIDTH                (512),
		.LENGTH_WIDTH              (20),
		.FIFO_DEPTH                (128),
		.STRIDE_ENABLE             (0),
		.BURST_ENABLE              (1),
		.PACKET_ENABLE             (0),
		.ERROR_ENABLE              (0),
		.ERROR_WIDTH               (8),
		.CHANNEL_ENABLE            (0),
		.CHANNEL_WIDTH             (8),
		.BYTE_ENABLE_WIDTH         (64),
		.BYTE_ENABLE_WIDTH_LOG2    (6),
		.ADDRESS_WIDTH             (34),
		.FIFO_DEPTH_LOG2           (7),
		.SYMBOL_WIDTH              (8),
		.NUMBER_OF_SYMBOLS         (64),
		.NUMBER_OF_SYMBOLS_LOG2    (6),
		.MAX_BURST_COUNT_WIDTH     (5),
		.UNALIGNED_ACCESSES_ENABLE (0),
		.ONLY_FULL_ACCESS_ENABLE   (1),
		.BURST_WRAPPING_SUPPORT    (1),
		.PROGRAMMABLE_BURST_ENABLE (0),
		.MAX_BURST_COUNT           (16),
		.FIFO_SPEED_OPTIMIZATION   (1),
		.STRIDE_WIDTH              (1)
	) dma_read_master (
		.clk                  (dma_clk_clk),                                          //            Clock.clk
		.reset                (~dma_reset_reset_n),                                   //      Clock_reset.reset
		.master_address       (dma_read_master_data_read_master_address),             // Data_Read_Master.address
		.master_read          (dma_read_master_data_read_master_read),                //                 .read
		.master_byteenable    (dma_read_master_data_read_master_byteenable),          //                 .byteenable
		.master_readdata      (dma_read_master_data_read_master_readdata),            //                 .readdata
		.master_waitrequest   (dma_read_master_data_read_master_waitrequest),         //                 .waitrequest
		.master_readdatavalid (dma_read_master_data_read_master_readdatavalid),       //                 .readdatavalid
		.master_burstcount    (dma_read_master_data_read_master_burstcount),          //                 .burstcount
		.src_data             (dma_read_master_data_source_data),                     //      Data_Source.data
		.src_valid            (dma_read_master_data_source_valid),                    //                 .valid
		.src_ready            (dma_read_master_data_source_ready),                    //                 .ready
		.snk_command_data     (modular_sgdma_dispatcher_0_read_command_source_data),  //     Command_Sink.data
		.snk_command_valid    (modular_sgdma_dispatcher_0_read_command_source_valid), //                 .valid
		.snk_command_ready    (modular_sgdma_dispatcher_0_read_command_source_ready), //                 .ready
		.src_response_data    (dma_read_master_response_source_data),                 //  Response_Source.data
		.src_response_valid   (dma_read_master_response_source_valid),                //                 .valid
		.src_response_ready   (dma_read_master_response_source_ready),                //                 .ready
		.src_sop              (),                                                     //      (terminated)
		.src_eop              (),                                                     //      (terminated)
		.src_empty            (),                                                     //      (terminated)
		.src_error            (),                                                     //      (terminated)
		.src_channel          ()                                                      //      (terminated)
	);

	write_master #(
		.DATA_WIDTH                     (512),
		.LENGTH_WIDTH                   (20),
		.FIFO_DEPTH                     (128),
		.STRIDE_ENABLE                  (0),
		.BURST_ENABLE                   (1),
		.PACKET_ENABLE                  (0),
		.ERROR_ENABLE                   (0),
		.ERROR_WIDTH                    (8),
		.BYTE_ENABLE_WIDTH              (64),
		.BYTE_ENABLE_WIDTH_LOG2         (6),
		.ADDRESS_WIDTH                  (34),
		.FIFO_DEPTH_LOG2                (7),
		.SYMBOL_WIDTH                   (8),
		.NUMBER_OF_SYMBOLS              (64),
		.NUMBER_OF_SYMBOLS_LOG2         (6),
		.MAX_BURST_COUNT_WIDTH          (5),
		.UNALIGNED_ACCESSES_ENABLE      (0),
		.ONLY_FULL_ACCESS_ENABLE        (1),
		.BURST_WRAPPING_SUPPORT         (1),
		.PROGRAMMABLE_BURST_ENABLE      (0),
		.MAX_BURST_COUNT                (16),
		.FIFO_SPEED_OPTIMIZATION        (1),
		.STRIDE_WIDTH                   (1),
		.ACTUAL_BYTES_TRANSFERRED_WIDTH (32)
	) dma_write_master (
		.clk                (dma_clk_clk),                                           //             Clock.clk
		.reset              (~dma_reset_reset_n),                                    //       Clock_reset.reset
		.master_address     (dma_write_master_data_write_master_address),            // Data_Write_Master.address
		.master_write       (dma_write_master_data_write_master_write),              //                  .write
		.master_byteenable  (dma_write_master_data_write_master_byteenable),         //                  .byteenable
		.master_writedata   (dma_write_master_data_write_master_writedata),          //                  .writedata
		.master_waitrequest (dma_write_master_data_write_master_waitrequest),        //                  .waitrequest
		.master_burstcount  (dma_write_master_data_write_master_burstcount),         //                  .burstcount
		.snk_data           (dma_read_master_data_source_data),                      //         Data_Sink.data
		.snk_valid          (dma_read_master_data_source_valid),                     //                  .valid
		.snk_ready          (dma_read_master_data_source_ready),                     //                  .ready
		.snk_command_data   (modular_sgdma_dispatcher_0_write_command_source_data),  //      Command_Sink.data
		.snk_command_valid  (modular_sgdma_dispatcher_0_write_command_source_valid), //                  .valid
		.snk_command_ready  (modular_sgdma_dispatcher_0_write_command_source_ready), //                  .ready
		.src_response_data  (dma_write_master_response_source_data),                 //   Response_Source.data
		.src_response_valid (dma_write_master_response_source_valid),                //                  .valid
		.src_response_ready (dma_write_master_response_source_ready),                //                  .ready
		.snk_sop            (1'b0),                                                  //       (terminated)
		.snk_eop            (1'b0),                                                  //       (terminated)
		.snk_empty          (6'b000000),                                             //       (terminated)
		.snk_error          (8'b00000000)                                            //       (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (512),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (34),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pipe_stage_dma_read (
		.clk              (dma_clk_clk),                                            //   clk.clk
		.reset            (~dma_reset_reset_n),                                     // reset.reset
		.s0_waitrequest   (mm_interconnect_1_pipe_stage_dma_read_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_pipe_stage_dma_read_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_pipe_stage_dma_read_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_pipe_stage_dma_read_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_pipe_stage_dma_read_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_pipe_stage_dma_read_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_pipe_stage_dma_read_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_pipe_stage_dma_read_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_pipe_stage_dma_read_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_pipe_stage_dma_read_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (dma_read_waitrequest),                                   //    m0.waitrequest
		.m0_readdata      (dma_read_readdata),                                      //      .readdata
		.m0_readdatavalid (dma_read_readdatavalid),                                 //      .readdatavalid
		.m0_burstcount    (dma_read_burstcount),                                    //      .burstcount
		.m0_writedata     (dma_read_writedata),                                     //      .writedata
		.m0_address       (dma_read_address),                                       //      .address
		.m0_write         (dma_read_write),                                         //      .write
		.m0_read          (dma_read_read),                                          //      .read
		.m0_byteenable    (dma_read_byteenable),                                    //      .byteenable
		.m0_debugaccess   (dma_read_debugaccess),                                   //      .debugaccess
		.s0_response      (),                                                       // (terminated)
		.m0_response      (2'b00)                                                   // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (512),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (34),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pipe_stage_dma_write (
		.clk              (dma_clk_clk),                                             //   clk.clk
		.reset            (~dma_reset_reset_n),                                      // reset.reset
		.s0_waitrequest   (mm_interconnect_0_pipe_stage_dma_write_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_pipe_stage_dma_write_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_pipe_stage_dma_write_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_pipe_stage_dma_write_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_pipe_stage_dma_write_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_pipe_stage_dma_write_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_pipe_stage_dma_write_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_pipe_stage_dma_write_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_pipe_stage_dma_write_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_pipe_stage_dma_write_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (dma_write_waitrequest),                                   //    m0.waitrequest
		.m0_readdata      (dma_write_readdata),                                      //      .readdata
		.m0_readdatavalid (dma_write_readdatavalid),                                 //      .readdatavalid
		.m0_burstcount    (dma_write_burstcount),                                    //      .burstcount
		.m0_writedata     (dma_write_writedata),                                     //      .writedata
		.m0_address       (dma_write_address),                                       //      .address
		.m0_write         (dma_write_write),                                         //      .write
		.m0_read          (dma_write_read),                                          //      .read
		.m0_byteenable    (dma_write_byteenable),                                    //      .byteenable
		.m0_debugaccess   (dma_write_debugaccess),                                   //      .debugaccess
		.s0_response      (),                                                        // (terminated)
		.m0_response      (2'b00)                                                    // (terminated)
	);

	system_acl_iface_dma_0_dma_mm_interconnect_0 mm_interconnect_0 (
		.dma_clk_clk_clk                                          (dma_clk_clk),                                             //                                        dma_clk_clk.clk
		.dma_write_master_Clock_reset_reset_bridge_in_reset_reset (~dma_reset_reset_n),                                      // dma_write_master_Clock_reset_reset_bridge_in_reset.reset
		.dma_write_master_Data_Write_Master_address               (dma_write_master_data_write_master_address),              //                 dma_write_master_Data_Write_Master.address
		.dma_write_master_Data_Write_Master_waitrequest           (dma_write_master_data_write_master_waitrequest),          //                                                   .waitrequest
		.dma_write_master_Data_Write_Master_burstcount            (dma_write_master_data_write_master_burstcount),           //                                                   .burstcount
		.dma_write_master_Data_Write_Master_byteenable            (dma_write_master_data_write_master_byteenable),           //                                                   .byteenable
		.dma_write_master_Data_Write_Master_write                 (dma_write_master_data_write_master_write),                //                                                   .write
		.dma_write_master_Data_Write_Master_writedata             (dma_write_master_data_write_master_writedata),            //                                                   .writedata
		.pipe_stage_dma_write_s0_address                          (mm_interconnect_0_pipe_stage_dma_write_s0_address),       //                            pipe_stage_dma_write_s0.address
		.pipe_stage_dma_write_s0_write                            (mm_interconnect_0_pipe_stage_dma_write_s0_write),         //                                                   .write
		.pipe_stage_dma_write_s0_read                             (mm_interconnect_0_pipe_stage_dma_write_s0_read),          //                                                   .read
		.pipe_stage_dma_write_s0_readdata                         (mm_interconnect_0_pipe_stage_dma_write_s0_readdata),      //                                                   .readdata
		.pipe_stage_dma_write_s0_writedata                        (mm_interconnect_0_pipe_stage_dma_write_s0_writedata),     //                                                   .writedata
		.pipe_stage_dma_write_s0_burstcount                       (mm_interconnect_0_pipe_stage_dma_write_s0_burstcount),    //                                                   .burstcount
		.pipe_stage_dma_write_s0_byteenable                       (mm_interconnect_0_pipe_stage_dma_write_s0_byteenable),    //                                                   .byteenable
		.pipe_stage_dma_write_s0_readdatavalid                    (mm_interconnect_0_pipe_stage_dma_write_s0_readdatavalid), //                                                   .readdatavalid
		.pipe_stage_dma_write_s0_waitrequest                      (mm_interconnect_0_pipe_stage_dma_write_s0_waitrequest),   //                                                   .waitrequest
		.pipe_stage_dma_write_s0_debugaccess                      (mm_interconnect_0_pipe_stage_dma_write_s0_debugaccess)    //                                                   .debugaccess
	);

	system_acl_iface_dma_0_dma_mm_interconnect_1 mm_interconnect_1 (
		.dma_clk_clk_clk                                         (dma_clk_clk),                                            //                                       dma_clk_clk.clk
		.dma_read_master_Clock_reset_reset_bridge_in_reset_reset (~dma_reset_reset_n),                                     // dma_read_master_Clock_reset_reset_bridge_in_reset.reset
		.dma_read_master_Data_Read_Master_address                (dma_read_master_data_read_master_address),               //                  dma_read_master_Data_Read_Master.address
		.dma_read_master_Data_Read_Master_waitrequest            (dma_read_master_data_read_master_waitrequest),           //                                                  .waitrequest
		.dma_read_master_Data_Read_Master_burstcount             (dma_read_master_data_read_master_burstcount),            //                                                  .burstcount
		.dma_read_master_Data_Read_Master_byteenable             (dma_read_master_data_read_master_byteenable),            //                                                  .byteenable
		.dma_read_master_Data_Read_Master_read                   (dma_read_master_data_read_master_read),                  //                                                  .read
		.dma_read_master_Data_Read_Master_readdata               (dma_read_master_data_read_master_readdata),              //                                                  .readdata
		.dma_read_master_Data_Read_Master_readdatavalid          (dma_read_master_data_read_master_readdatavalid),         //                                                  .readdatavalid
		.pipe_stage_dma_read_s0_address                          (mm_interconnect_1_pipe_stage_dma_read_s0_address),       //                            pipe_stage_dma_read_s0.address
		.pipe_stage_dma_read_s0_write                            (mm_interconnect_1_pipe_stage_dma_read_s0_write),         //                                                  .write
		.pipe_stage_dma_read_s0_read                             (mm_interconnect_1_pipe_stage_dma_read_s0_read),          //                                                  .read
		.pipe_stage_dma_read_s0_readdata                         (mm_interconnect_1_pipe_stage_dma_read_s0_readdata),      //                                                  .readdata
		.pipe_stage_dma_read_s0_writedata                        (mm_interconnect_1_pipe_stage_dma_read_s0_writedata),     //                                                  .writedata
		.pipe_stage_dma_read_s0_burstcount                       (mm_interconnect_1_pipe_stage_dma_read_s0_burstcount),    //                                                  .burstcount
		.pipe_stage_dma_read_s0_byteenable                       (mm_interconnect_1_pipe_stage_dma_read_s0_byteenable),    //                                                  .byteenable
		.pipe_stage_dma_read_s0_readdatavalid                    (mm_interconnect_1_pipe_stage_dma_read_s0_readdatavalid), //                                                  .readdatavalid
		.pipe_stage_dma_read_s0_waitrequest                      (mm_interconnect_1_pipe_stage_dma_read_s0_waitrequest),   //                                                  .waitrequest
		.pipe_stage_dma_read_s0_debugaccess                      (mm_interconnect_1_pipe_stage_dma_read_s0_debugaccess)    //                                                  .debugaccess
	);

endmodule

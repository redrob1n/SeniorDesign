// system_acl_iface.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module system_acl_iface (
		input  wire         reset_n,                               //               global_reset.reset_n
		input  wire         pcie_refclk_clk,                       //                pcie_refclk.clk
		input  wire         pcie_hip_serial_rx_in0,                //            pcie_hip_serial.rx_in0
		input  wire         pcie_hip_serial_rx_in1,                //                           .rx_in1
		input  wire         pcie_hip_serial_rx_in2,                //                           .rx_in2
		input  wire         pcie_hip_serial_rx_in3,                //                           .rx_in3
		input  wire         pcie_hip_serial_rx_in4,                //                           .rx_in4
		input  wire         pcie_hip_serial_rx_in5,                //                           .rx_in5
		input  wire         pcie_hip_serial_rx_in6,                //                           .rx_in6
		input  wire         pcie_hip_serial_rx_in7,                //                           .rx_in7
		output wire         pcie_hip_serial_tx_out0,               //                           .tx_out0
		output wire         pcie_hip_serial_tx_out1,               //                           .tx_out1
		output wire         pcie_hip_serial_tx_out2,               //                           .tx_out2
		output wire         pcie_hip_serial_tx_out3,               //                           .tx_out3
		output wire         pcie_hip_serial_tx_out4,               //                           .tx_out4
		output wire         pcie_hip_serial_tx_out5,               //                           .tx_out5
		output wire         pcie_hip_serial_tx_out6,               //                           .tx_out6
		output wire         pcie_hip_serial_tx_out7,               //                           .tx_out7
		input  wire         pcie_npor_npor,                        //                  pcie_npor.npor
		input  wire         pcie_npor_pin_perst,                   //                           .pin_perst
		output wire [14:0]  ddr3a_mem_a,                           //                      ddr3a.mem_a
		output wire [2:0]   ddr3a_mem_ba,                          //                           .mem_ba
		output wire [0:0]   ddr3a_mem_ck,                          //                           .mem_ck
		output wire [0:0]   ddr3a_mem_ck_n,                        //                           .mem_ck_n
		output wire [0:0]   ddr3a_mem_cke,                         //                           .mem_cke
		output wire [0:0]   ddr3a_mem_cs_n,                        //                           .mem_cs_n
		output wire [7:0]   ddr3a_mem_dm,                          //                           .mem_dm
		output wire [0:0]   ddr3a_mem_ras_n,                       //                           .mem_ras_n
		output wire [0:0]   ddr3a_mem_cas_n,                       //                           .mem_cas_n
		output wire [0:0]   ddr3a_mem_we_n,                        //                           .mem_we_n
		output wire         ddr3a_mem_reset_n,                     //                           .mem_reset_n
		inout  wire [63:0]  ddr3a_mem_dq,                          //                           .mem_dq
		inout  wire [7:0]   ddr3a_mem_dqs,                         //                           .mem_dqs
		inout  wire [7:0]   ddr3a_mem_dqs_n,                       //                           .mem_dqs_n
		output wire [0:0]   ddr3a_mem_odt,                         //                           .mem_odt
		input  wire         octa_rzqin,                            //                       octa.rzqin
		input  wire         ddr3a_pll_ref_clk,                     //              ddr3a_pll_ref.clk
		output wire [14:0]  ddr3b_mem_a,                           //                      ddr3b.mem_a
		output wire [2:0]   ddr3b_mem_ba,                          //                           .mem_ba
		output wire [0:0]   ddr3b_mem_ck,                          //                           .mem_ck
		output wire [0:0]   ddr3b_mem_ck_n,                        //                           .mem_ck_n
		output wire [0:0]   ddr3b_mem_cke,                         //                           .mem_cke
		output wire [0:0]   ddr3b_mem_cs_n,                        //                           .mem_cs_n
		output wire [7:0]   ddr3b_mem_dm,                          //                           .mem_dm
		output wire [0:0]   ddr3b_mem_ras_n,                       //                           .mem_ras_n
		output wire [0:0]   ddr3b_mem_cas_n,                       //                           .mem_cas_n
		output wire [0:0]   ddr3b_mem_we_n,                        //                           .mem_we_n
		output wire         ddr3b_mem_reset_n,                     //                           .mem_reset_n
		inout  wire [63:0]  ddr3b_mem_dq,                          //                           .mem_dq
		inout  wire [7:0]   ddr3b_mem_dqs,                         //                           .mem_dqs
		inout  wire [7:0]   ddr3b_mem_dqs_n,                       //                           .mem_dqs_n
		output wire [0:0]   ddr3b_mem_odt,                         //                           .mem_odt
		input  wire         octb_rzqin,                            //                       octb.rzqin
		input  wire         ddr3b_pll_ref_clk,                     //              ddr3b_pll_ref.clk
		input  wire [31:0]  pcie_hip_ctrl_test_in,                 //              pcie_hip_ctrl.test_in
		input  wire         pcie_hip_ctrl_simu_mode_pipe,          //                           .simu_mode_pipe
		input  wire         config_clk_clk,                        //                 config_clk.clk
		output wire [1:0]   acl_internal_memorg_kernel_mode,       // acl_internal_memorg_kernel.mode
		output wire         kernel_clk2x_clk,                      //               kernel_clk2x.clk
		input  wire         kernel_pll_refclk_clk,                 //          kernel_pll_refclk.clk
		input  wire         kernel_cra_waitrequest,                //                 kernel_cra.waitrequest
		input  wire [63:0]  kernel_cra_readdata,                   //                           .readdata
		input  wire         kernel_cra_readdatavalid,              //                           .readdatavalid
		output wire [0:0]   kernel_cra_burstcount,                 //                           .burstcount
		output wire [63:0]  kernel_cra_writedata,                  //                           .writedata
		output wire [29:0]  kernel_cra_address,                    //                           .address
		output wire         kernel_cra_write,                      //                           .write
		output wire         kernel_cra_read,                       //                           .read
		output wire [7:0]   kernel_cra_byteenable,                 //                           .byteenable
		output wire         kernel_cra_debugaccess,                //                           .debugaccess
		input  wire [0:0]   kernel_irq_irq,                        //                 kernel_irq.irq
		output wire         kernel_mem0_waitrequest,               //                kernel_mem0.waitrequest
		output wire [511:0] kernel_mem0_readdata,                  //                           .readdata
		output wire         kernel_mem0_readdatavalid,             //                           .readdatavalid
		input  wire [4:0]   kernel_mem0_burstcount,                //                           .burstcount
		input  wire [511:0] kernel_mem0_writedata,                 //                           .writedata
		input  wire [30:0]  kernel_mem0_address,                   //                           .address
		input  wire         kernel_mem0_write,                     //                           .write
		input  wire         kernel_mem0_read,                      //                           .read
		input  wire [63:0]  kernel_mem0_byteenable,                //                           .byteenable
		input  wire         kernel_mem0_debugaccess,               //                           .debugaccess
		output wire         kernel_mem1_waitrequest,               //                kernel_mem1.waitrequest
		output wire [511:0] kernel_mem1_readdata,                  //                           .readdata
		output wire         kernel_mem1_readdatavalid,             //                           .readdatavalid
		input  wire [4:0]   kernel_mem1_burstcount,                //                           .burstcount
		input  wire [511:0] kernel_mem1_writedata,                 //                           .writedata
		input  wire [30:0]  kernel_mem1_address,                   //                           .address
		input  wire         kernel_mem1_write,                     //                           .write
		input  wire         kernel_mem1_read,                      //                           .read
		input  wire [63:0]  kernel_mem1_byteenable,                //                           .byteenable
		input  wire         kernel_mem1_debugaccess,               //                           .debugaccess
		output wire [31:0]  acl_internal_snoop_data,               //         acl_internal_snoop.data
		output wire         acl_internal_snoop_valid,              //                           .valid
		input  wire         acl_internal_snoop_ready,              //                           .ready
		output wire         kernel_clk_clk,                        //                 kernel_clk.clk
		output wire         kernel_reset_reset_n,                  //               kernel_reset.reset_n
		output wire         pcie_npor_out_reset_n,                 //              pcie_npor_out.reset_n
		input  wire [699:0] reconfig_to_xcvr_reconfig_to_xcvr,     //           reconfig_to_xcvr.reconfig_to_xcvr
		output wire [459:0] reconfig_from_xcvr_reconfig_from_xcvr  //         reconfig_from_xcvr.reconfig_from_xcvr
	);

	wire          ddr3b_afi_clk_clk;                                                // ddr3b:afi_clk -> [clock_cross_dma_to_ddr3b:m0_clk, clock_cross_kernel_mem_1:m0_clk, em_pc_1:avl_clk, mm_interconnect_10:ddr3b_afi_clk_clk, mm_interconnect_1:ddr3b_afi_clk_clk, mm_interconnect_2:ddr3b_afi_clk_clk, mm_interconnect_7:ddr3b_afi_clk_clk, pipe_stage_ddr3b_dimm:clk, pipe_stage_ddr3b_iface:clk, reset_controller_ddr3b:clk, rst_controller_004:clk, rst_controller_007:clk]
	wire          ddr3a_afi_clk_clk;                                                // ddr3a:afi_clk -> [acl_memory_bank_divider_0:clk_clk, clock_cross_dma_to_ddr3b:s0_clk, clock_cross_dma_to_pcie:s0_clk, clock_cross_kernel_mem_0:m0_clk, dma_0:clk_clk, em_pc_0:avl_clk, irq_synchronizer_001:receiver_clk, mm_interconnect_0:ddr3a_afi_clk_clk, mm_interconnect_12:ddr3a_afi_clk_clk, mm_interconnect_2:ddr3a_afi_clk_clk, mm_interconnect_3:ddr3a_afi_clk_clk, mm_interconnect_5:ddr3a_afi_clk_clk, mm_interconnect_6:ddr3a_afi_clk_clk, pipe_stage_ddr3a_dimm:clk, pipe_stage_ddr3a_iface:clk, reset_controller_ddr3a:clk, rst_controller:clk, rst_controller_002:clk, rst_controller_003:clk]
	wire          pcie_coreclkout_clk;                                              // pcie:coreclkout -> [clock_cross_dma_to_pcie:m0_clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, kernel_interface:clk_clk, mm_interconnect_2:pcie_coreclkout_clk, mm_interconnect_8:pcie_coreclkout_clk, mm_interconnect_9:pcie_coreclkout_clk, pipe_stage_host_ctrl:clk, reset_controller_pcie:clk, rst_controller_006:clk, rst_controller_008:clk, uniphy_status_0:clk, version_id_0:clk]
	wire          temperature_pll_outclk0_clk;                                      // temperature_pll:outclk_0 -> [mm_interconnect_2:temperature_pll_outclk0_clk, rst_controller_001:clk, temperature_0:clk]
	wire          pipe_stage_ddr3a_iface_m0_waitrequest;                            // pipe_stage_ddr3a_dimm:s0_waitrequest -> pipe_stage_ddr3a_iface:m0_waitrequest
	wire  [511:0] pipe_stage_ddr3a_iface_m0_readdata;                               // pipe_stage_ddr3a_dimm:s0_readdata -> pipe_stage_ddr3a_iface:m0_readdata
	wire          pipe_stage_ddr3a_iface_m0_debugaccess;                            // pipe_stage_ddr3a_iface:m0_debugaccess -> pipe_stage_ddr3a_dimm:s0_debugaccess
	wire   [30:0] pipe_stage_ddr3a_iface_m0_address;                                // pipe_stage_ddr3a_iface:m0_address -> pipe_stage_ddr3a_dimm:s0_address
	wire          pipe_stage_ddr3a_iface_m0_read;                                   // pipe_stage_ddr3a_iface:m0_read -> pipe_stage_ddr3a_dimm:s0_read
	wire   [63:0] pipe_stage_ddr3a_iface_m0_byteenable;                             // pipe_stage_ddr3a_iface:m0_byteenable -> pipe_stage_ddr3a_dimm:s0_byteenable
	wire          pipe_stage_ddr3a_iface_m0_readdatavalid;                          // pipe_stage_ddr3a_dimm:s0_readdatavalid -> pipe_stage_ddr3a_iface:m0_readdatavalid
	wire  [511:0] pipe_stage_ddr3a_iface_m0_writedata;                              // pipe_stage_ddr3a_iface:m0_writedata -> pipe_stage_ddr3a_dimm:s0_writedata
	wire          pipe_stage_ddr3a_iface_m0_write;                                  // pipe_stage_ddr3a_iface:m0_write -> pipe_stage_ddr3a_dimm:s0_write
	wire    [4:0] pipe_stage_ddr3a_iface_m0_burstcount;                             // pipe_stage_ddr3a_iface:m0_burstcount -> pipe_stage_ddr3a_dimm:s0_burstcount
	wire    [1:0] kernel_interface_acl_bsp_memorg_host_mode;                        // kernel_interface:acl_bsp_memorg_host_mode -> acl_memory_bank_divider_0:acl_bsp_memorg_host_mode
	wire          reset_controller_pcie_reset_out_reset;                            // reset_controller_pcie:reset_out -> [clock_cross_dma_to_pcie:m0_reset, kernel_interface:reset_reset_n, kernel_interface:sw_reset_in_reset, mm_interconnect_2:pipe_stage_host_ctrl_reset_reset_bridge_in_reset_reset, mm_interconnect_8:pipe_stage_host_ctrl_reset_reset_bridge_in_reset_reset, mm_interconnect_9:clock_cross_dma_to_pcie_m0_reset_reset_bridge_in_reset_reset, pipe_stage_host_ctrl:reset, rst_controller_009:reset_in0]
	wire          reset_controller_ddr3a_reset_out_reset;                           // reset_controller_ddr3a:reset_out -> [clock_cross_dma_to_ddr3b:s0_reset, em_pc_0:avl_reset_n, mm_interconnect_0:pipe_stage_ddr3a_dimm_reset_reset_bridge_in_reset_reset, mm_interconnect_12:clock_cross_dma_to_ddr3b_s0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:em_pc_0_avl_reset_n_reset_bridge_in_reset_reset, mm_interconnect_2:em_pc_0_em_csr_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_5:em_pc_0_avl_in_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_5:em_pc_0_avl_reset_n_reset_bridge_in_reset_reset, mm_interconnect_6:em_pc_0_avl_reset_n_reset_bridge_in_reset_reset, mm_interconnect_6:pipe_stage_ddr3a_iface_reset_reset_bridge_in_reset_reset, pipe_stage_ddr3a_dimm:reset, pipe_stage_ddr3a_iface:reset]
	wire          reset_controller_ddr3b_reset_out_reset;                           // reset_controller_ddr3b:reset_out -> [clock_cross_dma_to_ddr3b:m0_reset, em_pc_1:avl_reset_n, mm_interconnect_10:clock_cross_dma_to_ddr3b_m0_reset_reset_bridge_in_reset_reset, mm_interconnect_10:em_pc_1_avl_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:pipe_stage_ddr3b_dimm_reset_reset_bridge_in_reset_reset, mm_interconnect_2:em_pc_1_avl_reset_n_reset_bridge_in_reset_reset, mm_interconnect_2:em_pc_1_em_csr_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_7:em_pc_1_avl_in_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_7:em_pc_1_avl_reset_n_reset_bridge_in_reset_reset, pipe_stage_ddr3b_dimm:reset, pipe_stage_ddr3b_iface:reset, rst_controller_002:reset_in0]
	wire          pcie_nreset_status_reset;                                         // pcie:reset_status -> [reset_controller_global:reset_in1, rst_controller_008:reset_in0]
	wire          reset_controller_global_reset_out_reset;                          // reset_controller_global:reset_out -> [acl_kernel_clk:reset_reset_n, ddr3a:global_reset_n, ddr3a:soft_reset_n, ddr3b:global_reset_n, ddr3b:soft_reset_n, mm_interconnect_2:acl_kernel_clk_reset_reset_bridge_in_reset_reset, reset_controller_ddr3a:reset_in0, reset_controller_ddr3b:reset_in0, reset_controller_pcie:reset_in0, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_006:reset_in0, rst_controller_007:reset_in0, temperature_pll:rst]
	wire          ddr3a_status_local_cal_fail;                                      // ddr3a:local_cal_fail -> uniphy_status_0:mem0_local_cal_fail
	wire          ddr3a_status_local_init_done;                                     // ddr3a:local_init_done -> uniphy_status_0:mem0_local_init_done
	wire          ddr3a_status_local_cal_success;                                   // ddr3a:local_cal_success -> uniphy_status_0:mem0_local_cal_success
	wire          ddr3b_status_local_cal_fail;                                      // ddr3b:local_cal_fail -> uniphy_status_0:mem1_local_cal_fail
	wire          ddr3b_status_local_init_done;                                     // ddr3b:local_init_done -> uniphy_status_0:mem1_local_init_done
	wire          ddr3b_status_local_cal_success;                                   // ddr3b:local_cal_success -> uniphy_status_0:mem1_local_cal_success
	wire          pipe_stage_ddr3b_iface_m0_waitrequest;                            // pipe_stage_ddr3b_dimm:s0_waitrequest -> pipe_stage_ddr3b_iface:m0_waitrequest
	wire  [511:0] pipe_stage_ddr3b_iface_m0_readdata;                               // pipe_stage_ddr3b_dimm:s0_readdata -> pipe_stage_ddr3b_iface:m0_readdata
	wire          pipe_stage_ddr3b_iface_m0_debugaccess;                            // pipe_stage_ddr3b_iface:m0_debugaccess -> pipe_stage_ddr3b_dimm:s0_debugaccess
	wire   [30:0] pipe_stage_ddr3b_iface_m0_address;                                // pipe_stage_ddr3b_iface:m0_address -> pipe_stage_ddr3b_dimm:s0_address
	wire          pipe_stage_ddr3b_iface_m0_read;                                   // pipe_stage_ddr3b_iface:m0_read -> pipe_stage_ddr3b_dimm:s0_read
	wire   [63:0] pipe_stage_ddr3b_iface_m0_byteenable;                             // pipe_stage_ddr3b_iface:m0_byteenable -> pipe_stage_ddr3b_dimm:s0_byteenable
	wire          pipe_stage_ddr3b_iface_m0_readdatavalid;                          // pipe_stage_ddr3b_dimm:s0_readdatavalid -> pipe_stage_ddr3b_iface:m0_readdatavalid
	wire  [511:0] pipe_stage_ddr3b_iface_m0_writedata;                              // pipe_stage_ddr3b_iface:m0_writedata -> pipe_stage_ddr3b_dimm:s0_writedata
	wire          pipe_stage_ddr3b_iface_m0_write;                                  // pipe_stage_ddr3b_iface:m0_write -> pipe_stage_ddr3b_dimm:s0_write
	wire    [4:0] pipe_stage_ddr3b_iface_m0_burstcount;                             // pipe_stage_ddr3b_iface:m0_burstcount -> pipe_stage_ddr3b_dimm:s0_burstcount
	wire          pipe_stage_ddr3a_dimm_m0_waitrequest;                             // mm_interconnect_0:pipe_stage_ddr3a_dimm_m0_waitrequest -> pipe_stage_ddr3a_dimm:m0_waitrequest
	wire  [511:0] pipe_stage_ddr3a_dimm_m0_readdata;                                // mm_interconnect_0:pipe_stage_ddr3a_dimm_m0_readdata -> pipe_stage_ddr3a_dimm:m0_readdata
	wire          pipe_stage_ddr3a_dimm_m0_debugaccess;                             // pipe_stage_ddr3a_dimm:m0_debugaccess -> mm_interconnect_0:pipe_stage_ddr3a_dimm_m0_debugaccess
	wire   [30:0] pipe_stage_ddr3a_dimm_m0_address;                                 // pipe_stage_ddr3a_dimm:m0_address -> mm_interconnect_0:pipe_stage_ddr3a_dimm_m0_address
	wire          pipe_stage_ddr3a_dimm_m0_read;                                    // pipe_stage_ddr3a_dimm:m0_read -> mm_interconnect_0:pipe_stage_ddr3a_dimm_m0_read
	wire   [63:0] pipe_stage_ddr3a_dimm_m0_byteenable;                              // pipe_stage_ddr3a_dimm:m0_byteenable -> mm_interconnect_0:pipe_stage_ddr3a_dimm_m0_byteenable
	wire          pipe_stage_ddr3a_dimm_m0_readdatavalid;                           // mm_interconnect_0:pipe_stage_ddr3a_dimm_m0_readdatavalid -> pipe_stage_ddr3a_dimm:m0_readdatavalid
	wire  [511:0] pipe_stage_ddr3a_dimm_m0_writedata;                               // pipe_stage_ddr3a_dimm:m0_writedata -> mm_interconnect_0:pipe_stage_ddr3a_dimm_m0_writedata
	wire          pipe_stage_ddr3a_dimm_m0_write;                                   // pipe_stage_ddr3a_dimm:m0_write -> mm_interconnect_0:pipe_stage_ddr3a_dimm_m0_write
	wire    [4:0] pipe_stage_ddr3a_dimm_m0_burstcount;                              // pipe_stage_ddr3a_dimm:m0_burstcount -> mm_interconnect_0:pipe_stage_ddr3a_dimm_m0_burstcount
	wire          mm_interconnect_0_ddr3a_avl_beginbursttransfer;                   // mm_interconnect_0:ddr3a_avl_beginbursttransfer -> ddr3a:avl_burstbegin
	wire  [511:0] mm_interconnect_0_ddr3a_avl_readdata;                             // ddr3a:avl_rdata -> mm_interconnect_0:ddr3a_avl_readdata
	wire          mm_interconnect_0_ddr3a_avl_waitrequest;                          // ddr3a:avl_ready -> mm_interconnect_0:ddr3a_avl_waitrequest
	wire   [24:0] mm_interconnect_0_ddr3a_avl_address;                              // mm_interconnect_0:ddr3a_avl_address -> ddr3a:avl_addr
	wire          mm_interconnect_0_ddr3a_avl_read;                                 // mm_interconnect_0:ddr3a_avl_read -> ddr3a:avl_read_req
	wire   [63:0] mm_interconnect_0_ddr3a_avl_byteenable;                           // mm_interconnect_0:ddr3a_avl_byteenable -> ddr3a:avl_be
	wire          mm_interconnect_0_ddr3a_avl_readdatavalid;                        // ddr3a:avl_rdata_valid -> mm_interconnect_0:ddr3a_avl_readdatavalid
	wire          mm_interconnect_0_ddr3a_avl_write;                                // mm_interconnect_0:ddr3a_avl_write -> ddr3a:avl_write_req
	wire  [511:0] mm_interconnect_0_ddr3a_avl_writedata;                            // mm_interconnect_0:ddr3a_avl_writedata -> ddr3a:avl_wdata
	wire    [4:0] mm_interconnect_0_ddr3a_avl_burstcount;                           // mm_interconnect_0:ddr3a_avl_burstcount -> ddr3a:avl_size
	wire          pipe_stage_ddr3b_dimm_m0_waitrequest;                             // mm_interconnect_1:pipe_stage_ddr3b_dimm_m0_waitrequest -> pipe_stage_ddr3b_dimm:m0_waitrequest
	wire  [511:0] pipe_stage_ddr3b_dimm_m0_readdata;                                // mm_interconnect_1:pipe_stage_ddr3b_dimm_m0_readdata -> pipe_stage_ddr3b_dimm:m0_readdata
	wire          pipe_stage_ddr3b_dimm_m0_debugaccess;                             // pipe_stage_ddr3b_dimm:m0_debugaccess -> mm_interconnect_1:pipe_stage_ddr3b_dimm_m0_debugaccess
	wire   [30:0] pipe_stage_ddr3b_dimm_m0_address;                                 // pipe_stage_ddr3b_dimm:m0_address -> mm_interconnect_1:pipe_stage_ddr3b_dimm_m0_address
	wire          pipe_stage_ddr3b_dimm_m0_read;                                    // pipe_stage_ddr3b_dimm:m0_read -> mm_interconnect_1:pipe_stage_ddr3b_dimm_m0_read
	wire   [63:0] pipe_stage_ddr3b_dimm_m0_byteenable;                              // pipe_stage_ddr3b_dimm:m0_byteenable -> mm_interconnect_1:pipe_stage_ddr3b_dimm_m0_byteenable
	wire          pipe_stage_ddr3b_dimm_m0_readdatavalid;                           // mm_interconnect_1:pipe_stage_ddr3b_dimm_m0_readdatavalid -> pipe_stage_ddr3b_dimm:m0_readdatavalid
	wire  [511:0] pipe_stage_ddr3b_dimm_m0_writedata;                               // pipe_stage_ddr3b_dimm:m0_writedata -> mm_interconnect_1:pipe_stage_ddr3b_dimm_m0_writedata
	wire          pipe_stage_ddr3b_dimm_m0_write;                                   // pipe_stage_ddr3b_dimm:m0_write -> mm_interconnect_1:pipe_stage_ddr3b_dimm_m0_write
	wire    [4:0] pipe_stage_ddr3b_dimm_m0_burstcount;                              // pipe_stage_ddr3b_dimm:m0_burstcount -> mm_interconnect_1:pipe_stage_ddr3b_dimm_m0_burstcount
	wire          mm_interconnect_1_ddr3b_avl_beginbursttransfer;                   // mm_interconnect_1:ddr3b_avl_beginbursttransfer -> ddr3b:avl_burstbegin
	wire  [511:0] mm_interconnect_1_ddr3b_avl_readdata;                             // ddr3b:avl_rdata -> mm_interconnect_1:ddr3b_avl_readdata
	wire          mm_interconnect_1_ddr3b_avl_waitrequest;                          // ddr3b:avl_ready -> mm_interconnect_1:ddr3b_avl_waitrequest
	wire   [24:0] mm_interconnect_1_ddr3b_avl_address;                              // mm_interconnect_1:ddr3b_avl_address -> ddr3b:avl_addr
	wire          mm_interconnect_1_ddr3b_avl_read;                                 // mm_interconnect_1:ddr3b_avl_read -> ddr3b:avl_read_req
	wire   [63:0] mm_interconnect_1_ddr3b_avl_byteenable;                           // mm_interconnect_1:ddr3b_avl_byteenable -> ddr3b:avl_be
	wire          mm_interconnect_1_ddr3b_avl_readdatavalid;                        // ddr3b:avl_rdata_valid -> mm_interconnect_1:ddr3b_avl_readdatavalid
	wire          mm_interconnect_1_ddr3b_avl_write;                                // mm_interconnect_1:ddr3b_avl_write -> ddr3b:avl_write_req
	wire  [511:0] mm_interconnect_1_ddr3b_avl_writedata;                            // mm_interconnect_1:ddr3b_avl_writedata -> ddr3b:avl_wdata
	wire    [4:0] mm_interconnect_1_ddr3b_avl_burstcount;                           // mm_interconnect_1:ddr3b_avl_burstcount -> ddr3b:avl_size
	wire          pipe_stage_host_ctrl_m0_waitrequest;                              // mm_interconnect_2:pipe_stage_host_ctrl_m0_waitrequest -> pipe_stage_host_ctrl:m0_waitrequest
	wire   [31:0] pipe_stage_host_ctrl_m0_readdata;                                 // mm_interconnect_2:pipe_stage_host_ctrl_m0_readdata -> pipe_stage_host_ctrl:m0_readdata
	wire          pipe_stage_host_ctrl_m0_debugaccess;                              // pipe_stage_host_ctrl:m0_debugaccess -> mm_interconnect_2:pipe_stage_host_ctrl_m0_debugaccess
	wire   [17:0] pipe_stage_host_ctrl_m0_address;                                  // pipe_stage_host_ctrl:m0_address -> mm_interconnect_2:pipe_stage_host_ctrl_m0_address
	wire          pipe_stage_host_ctrl_m0_read;                                     // pipe_stage_host_ctrl:m0_read -> mm_interconnect_2:pipe_stage_host_ctrl_m0_read
	wire    [3:0] pipe_stage_host_ctrl_m0_byteenable;                               // pipe_stage_host_ctrl:m0_byteenable -> mm_interconnect_2:pipe_stage_host_ctrl_m0_byteenable
	wire          pipe_stage_host_ctrl_m0_readdatavalid;                            // mm_interconnect_2:pipe_stage_host_ctrl_m0_readdatavalid -> pipe_stage_host_ctrl:m0_readdatavalid
	wire   [31:0] pipe_stage_host_ctrl_m0_writedata;                                // pipe_stage_host_ctrl:m0_writedata -> mm_interconnect_2:pipe_stage_host_ctrl_m0_writedata
	wire          pipe_stage_host_ctrl_m0_write;                                    // pipe_stage_host_ctrl:m0_write -> mm_interconnect_2:pipe_stage_host_ctrl_m0_write
	wire    [0:0] pipe_stage_host_ctrl_m0_burstcount;                               // pipe_stage_host_ctrl:m0_burstcount -> mm_interconnect_2:pipe_stage_host_ctrl_m0_burstcount
	wire   [31:0] mm_interconnect_2_temperature_0_s_readdata;                       // temperature_0:slave_readdata -> mm_interconnect_2:temperature_0_s_readdata
	wire          mm_interconnect_2_temperature_0_s_waitrequest;                    // temperature_0:slave_waitrequest -> mm_interconnect_2:temperature_0_s_waitrequest
	wire    [0:0] mm_interconnect_2_temperature_0_s_address;                        // mm_interconnect_2:temperature_0_s_address -> temperature_0:slave_address
	wire          mm_interconnect_2_temperature_0_s_read;                           // mm_interconnect_2:temperature_0_s_read -> temperature_0:slave_read
	wire    [3:0] mm_interconnect_2_temperature_0_s_byteenable;                     // mm_interconnect_2:temperature_0_s_byteenable -> temperature_0:slave_byteenable
	wire          mm_interconnect_2_temperature_0_s_readdatavalid;                  // temperature_0:slave_readdatavalid -> mm_interconnect_2:temperature_0_s_readdatavalid
	wire          mm_interconnect_2_temperature_0_s_write;                          // mm_interconnect_2:temperature_0_s_write -> temperature_0:slave_write
	wire   [31:0] mm_interconnect_2_temperature_0_s_writedata;                      // mm_interconnect_2:temperature_0_s_writedata -> temperature_0:slave_writedata
	wire   [31:0] mm_interconnect_2_acl_kernel_clk_ctrl_readdata;                   // acl_kernel_clk:ctrl_readdata -> mm_interconnect_2:acl_kernel_clk_ctrl_readdata
	wire          mm_interconnect_2_acl_kernel_clk_ctrl_waitrequest;                // acl_kernel_clk:ctrl_waitrequest -> mm_interconnect_2:acl_kernel_clk_ctrl_waitrequest
	wire          mm_interconnect_2_acl_kernel_clk_ctrl_debugaccess;                // mm_interconnect_2:acl_kernel_clk_ctrl_debugaccess -> acl_kernel_clk:ctrl_debugaccess
	wire   [10:0] mm_interconnect_2_acl_kernel_clk_ctrl_address;                    // mm_interconnect_2:acl_kernel_clk_ctrl_address -> acl_kernel_clk:ctrl_address
	wire          mm_interconnect_2_acl_kernel_clk_ctrl_read;                       // mm_interconnect_2:acl_kernel_clk_ctrl_read -> acl_kernel_clk:ctrl_read
	wire    [3:0] mm_interconnect_2_acl_kernel_clk_ctrl_byteenable;                 // mm_interconnect_2:acl_kernel_clk_ctrl_byteenable -> acl_kernel_clk:ctrl_byteenable
	wire          mm_interconnect_2_acl_kernel_clk_ctrl_readdatavalid;              // acl_kernel_clk:ctrl_readdatavalid -> mm_interconnect_2:acl_kernel_clk_ctrl_readdatavalid
	wire          mm_interconnect_2_acl_kernel_clk_ctrl_write;                      // mm_interconnect_2:acl_kernel_clk_ctrl_write -> acl_kernel_clk:ctrl_write
	wire   [31:0] mm_interconnect_2_acl_kernel_clk_ctrl_writedata;                  // mm_interconnect_2:acl_kernel_clk_ctrl_writedata -> acl_kernel_clk:ctrl_writedata
	wire    [0:0] mm_interconnect_2_acl_kernel_clk_ctrl_burstcount;                 // mm_interconnect_2:acl_kernel_clk_ctrl_burstcount -> acl_kernel_clk:ctrl_burstcount
	wire   [31:0] mm_interconnect_2_kernel_interface_kernel_cntrl_readdata;         // kernel_interface:kernel_cntrl_readdata -> mm_interconnect_2:kernel_interface_kernel_cntrl_readdata
	wire          mm_interconnect_2_kernel_interface_kernel_cntrl_waitrequest;      // kernel_interface:kernel_cntrl_waitrequest -> mm_interconnect_2:kernel_interface_kernel_cntrl_waitrequest
	wire          mm_interconnect_2_kernel_interface_kernel_cntrl_debugaccess;      // mm_interconnect_2:kernel_interface_kernel_cntrl_debugaccess -> kernel_interface:kernel_cntrl_debugaccess
	wire   [13:0] mm_interconnect_2_kernel_interface_kernel_cntrl_address;          // mm_interconnect_2:kernel_interface_kernel_cntrl_address -> kernel_interface:kernel_cntrl_address
	wire          mm_interconnect_2_kernel_interface_kernel_cntrl_read;             // mm_interconnect_2:kernel_interface_kernel_cntrl_read -> kernel_interface:kernel_cntrl_read
	wire    [3:0] mm_interconnect_2_kernel_interface_kernel_cntrl_byteenable;       // mm_interconnect_2:kernel_interface_kernel_cntrl_byteenable -> kernel_interface:kernel_cntrl_byteenable
	wire          mm_interconnect_2_kernel_interface_kernel_cntrl_readdatavalid;    // kernel_interface:kernel_cntrl_readdatavalid -> mm_interconnect_2:kernel_interface_kernel_cntrl_readdatavalid
	wire          mm_interconnect_2_kernel_interface_kernel_cntrl_write;            // mm_interconnect_2:kernel_interface_kernel_cntrl_write -> kernel_interface:kernel_cntrl_write
	wire   [31:0] mm_interconnect_2_kernel_interface_kernel_cntrl_writedata;        // mm_interconnect_2:kernel_interface_kernel_cntrl_writedata -> kernel_interface:kernel_cntrl_writedata
	wire    [0:0] mm_interconnect_2_kernel_interface_kernel_cntrl_burstcount;       // mm_interconnect_2:kernel_interface_kernel_cntrl_burstcount -> kernel_interface:kernel_cntrl_burstcount
	wire   [63:0] mm_interconnect_2_dma_0_csr_readdata;                             // dma_0:csr_readdata -> mm_interconnect_2:dma_0_csr_readdata
	wire          mm_interconnect_2_dma_0_csr_waitrequest;                          // dma_0:csr_waitrequest -> mm_interconnect_2:dma_0_csr_waitrequest
	wire          mm_interconnect_2_dma_0_csr_debugaccess;                          // mm_interconnect_2:dma_0_csr_debugaccess -> dma_0:csr_debugaccess
	wire    [9:0] mm_interconnect_2_dma_0_csr_address;                              // mm_interconnect_2:dma_0_csr_address -> dma_0:csr_address
	wire          mm_interconnect_2_dma_0_csr_read;                                 // mm_interconnect_2:dma_0_csr_read -> dma_0:csr_read
	wire    [7:0] mm_interconnect_2_dma_0_csr_byteenable;                           // mm_interconnect_2:dma_0_csr_byteenable -> dma_0:csr_byteenable
	wire          mm_interconnect_2_dma_0_csr_readdatavalid;                        // dma_0:csr_readdatavalid -> mm_interconnect_2:dma_0_csr_readdatavalid
	wire          mm_interconnect_2_dma_0_csr_write;                                // mm_interconnect_2:dma_0_csr_write -> dma_0:csr_write
	wire   [63:0] mm_interconnect_2_dma_0_csr_writedata;                            // mm_interconnect_2:dma_0_csr_writedata -> dma_0:csr_writedata
	wire    [0:0] mm_interconnect_2_dma_0_csr_burstcount;                           // mm_interconnect_2:dma_0_csr_burstcount -> dma_0:csr_burstcount
	wire          mm_interconnect_2_pcie_cra_chipselect;                            // mm_interconnect_2:pcie_Cra_chipselect -> pcie:CraChipSelect_i
	wire   [31:0] mm_interconnect_2_pcie_cra_readdata;                              // pcie:CraReadData_o -> mm_interconnect_2:pcie_Cra_readdata
	wire          mm_interconnect_2_pcie_cra_waitrequest;                           // pcie:CraWaitRequest_o -> mm_interconnect_2:pcie_Cra_waitrequest
	wire   [13:0] mm_interconnect_2_pcie_cra_address;                               // mm_interconnect_2:pcie_Cra_address -> pcie:CraAddress_i
	wire          mm_interconnect_2_pcie_cra_read;                                  // mm_interconnect_2:pcie_Cra_read -> pcie:CraRead
	wire    [3:0] mm_interconnect_2_pcie_cra_byteenable;                            // mm_interconnect_2:pcie_Cra_byteenable -> pcie:CraByteEnable_i
	wire          mm_interconnect_2_pcie_cra_write;                                 // mm_interconnect_2:pcie_Cra_write -> pcie:CraWrite
	wire   [31:0] mm_interconnect_2_pcie_cra_writedata;                             // mm_interconnect_2:pcie_Cra_writedata -> pcie:CraWriteData_i
	wire   [31:0] mm_interconnect_2_em_pc_0_em_csr_readdata;                        // em_pc_0:em_csr_readdata -> mm_interconnect_2:em_pc_0_em_csr_readdata
	wire          mm_interconnect_2_em_pc_0_em_csr_waitrequest;                     // em_pc_0:em_csr_waitrequest -> mm_interconnect_2:em_pc_0_em_csr_waitrequest
	wire          mm_interconnect_2_em_pc_0_em_csr_debugaccess;                     // mm_interconnect_2:em_pc_0_em_csr_debugaccess -> em_pc_0:em_csr_debugaccess
	wire   [13:0] mm_interconnect_2_em_pc_0_em_csr_address;                         // mm_interconnect_2:em_pc_0_em_csr_address -> em_pc_0:em_csr_address
	wire          mm_interconnect_2_em_pc_0_em_csr_read;                            // mm_interconnect_2:em_pc_0_em_csr_read -> em_pc_0:em_csr_read
	wire    [3:0] mm_interconnect_2_em_pc_0_em_csr_byteenable;                      // mm_interconnect_2:em_pc_0_em_csr_byteenable -> em_pc_0:em_csr_byteenable
	wire          mm_interconnect_2_em_pc_0_em_csr_readdatavalid;                   // em_pc_0:em_csr_readdatavalid -> mm_interconnect_2:em_pc_0_em_csr_readdatavalid
	wire          mm_interconnect_2_em_pc_0_em_csr_write;                           // mm_interconnect_2:em_pc_0_em_csr_write -> em_pc_0:em_csr_write
	wire   [31:0] mm_interconnect_2_em_pc_0_em_csr_writedata;                       // mm_interconnect_2:em_pc_0_em_csr_writedata -> em_pc_0:em_csr_writedata
	wire    [0:0] mm_interconnect_2_em_pc_0_em_csr_burstcount;                      // mm_interconnect_2:em_pc_0_em_csr_burstcount -> em_pc_0:em_csr_burstcount
	wire   [31:0] mm_interconnect_2_em_pc_1_em_csr_readdata;                        // em_pc_1:em_csr_readdata -> mm_interconnect_2:em_pc_1_em_csr_readdata
	wire          mm_interconnect_2_em_pc_1_em_csr_waitrequest;                     // em_pc_1:em_csr_waitrequest -> mm_interconnect_2:em_pc_1_em_csr_waitrequest
	wire          mm_interconnect_2_em_pc_1_em_csr_debugaccess;                     // mm_interconnect_2:em_pc_1_em_csr_debugaccess -> em_pc_1:em_csr_debugaccess
	wire   [13:0] mm_interconnect_2_em_pc_1_em_csr_address;                         // mm_interconnect_2:em_pc_1_em_csr_address -> em_pc_1:em_csr_address
	wire          mm_interconnect_2_em_pc_1_em_csr_read;                            // mm_interconnect_2:em_pc_1_em_csr_read -> em_pc_1:em_csr_read
	wire    [3:0] mm_interconnect_2_em_pc_1_em_csr_byteenable;                      // mm_interconnect_2:em_pc_1_em_csr_byteenable -> em_pc_1:em_csr_byteenable
	wire          mm_interconnect_2_em_pc_1_em_csr_readdatavalid;                   // em_pc_1:em_csr_readdatavalid -> mm_interconnect_2:em_pc_1_em_csr_readdatavalid
	wire          mm_interconnect_2_em_pc_1_em_csr_write;                           // mm_interconnect_2:em_pc_1_em_csr_write -> em_pc_1:em_csr_write
	wire   [31:0] mm_interconnect_2_em_pc_1_em_csr_writedata;                       // mm_interconnect_2:em_pc_1_em_csr_writedata -> em_pc_1:em_csr_writedata
	wire    [0:0] mm_interconnect_2_em_pc_1_em_csr_burstcount;                      // mm_interconnect_2:em_pc_1_em_csr_burstcount -> em_pc_1:em_csr_burstcount
	wire  [511:0] mm_interconnect_2_dma_0_s_nondma_readdata;                        // dma_0:s_nondma_readdata -> mm_interconnect_2:dma_0_s_nondma_readdata
	wire          mm_interconnect_2_dma_0_s_nondma_waitrequest;                     // dma_0:s_nondma_waitrequest -> mm_interconnect_2:dma_0_s_nondma_waitrequest
	wire    [9:0] mm_interconnect_2_dma_0_s_nondma_address;                         // mm_interconnect_2:dma_0_s_nondma_address -> dma_0:s_nondma_address
	wire          mm_interconnect_2_dma_0_s_nondma_read;                            // mm_interconnect_2:dma_0_s_nondma_read -> dma_0:s_nondma_read
	wire   [63:0] mm_interconnect_2_dma_0_s_nondma_byteenable;                      // mm_interconnect_2:dma_0_s_nondma_byteenable -> dma_0:s_nondma_byteenable
	wire          mm_interconnect_2_dma_0_s_nondma_readdatavalid;                   // dma_0:s_nondma_readdatavalid -> mm_interconnect_2:dma_0_s_nondma_readdatavalid
	wire          mm_interconnect_2_dma_0_s_nondma_write;                           // mm_interconnect_2:dma_0_s_nondma_write -> dma_0:s_nondma_write
	wire  [511:0] mm_interconnect_2_dma_0_s_nondma_writedata;                       // mm_interconnect_2:dma_0_s_nondma_writedata -> dma_0:s_nondma_writedata
	wire    [4:0] mm_interconnect_2_dma_0_s_nondma_burstcount;                      // mm_interconnect_2:dma_0_s_nondma_burstcount -> dma_0:s_nondma_burstcount
	wire   [31:0] mm_interconnect_2_uniphy_status_0_s_readdata;                     // uniphy_status_0:slave_readdata -> mm_interconnect_2:uniphy_status_0_s_readdata
	wire          mm_interconnect_2_uniphy_status_0_s_read;                         // mm_interconnect_2:uniphy_status_0_s_read -> uniphy_status_0:slave_read
	wire   [31:0] mm_interconnect_2_version_id_0_s_readdata;                        // version_id_0:slave_readdata -> mm_interconnect_2:version_id_0_s_readdata
	wire          mm_interconnect_2_version_id_0_s_read;                            // mm_interconnect_2:version_id_0_s_read -> version_id_0:slave_read
	wire          dma_0_m_waitrequest;                                              // mm_interconnect_3:dma_0_m_waitrequest -> dma_0:m_waitrequest
	wire  [511:0] dma_0_m_readdata;                                                 // mm_interconnect_3:dma_0_m_readdata -> dma_0:m_readdata
	wire          dma_0_m_debugaccess;                                              // dma_0:m_debugaccess -> mm_interconnect_3:dma_0_m_debugaccess
	wire   [33:0] dma_0_m_address;                                                  // dma_0:m_address -> mm_interconnect_3:dma_0_m_address
	wire          dma_0_m_read;                                                     // dma_0:m_read -> mm_interconnect_3:dma_0_m_read
	wire   [63:0] dma_0_m_byteenable;                                               // dma_0:m_byteenable -> mm_interconnect_3:dma_0_m_byteenable
	wire          dma_0_m_readdatavalid;                                            // mm_interconnect_3:dma_0_m_readdatavalid -> dma_0:m_readdatavalid
	wire  [511:0] dma_0_m_writedata;                                                // dma_0:m_writedata -> mm_interconnect_3:dma_0_m_writedata
	wire          dma_0_m_write;                                                    // dma_0:m_write -> mm_interconnect_3:dma_0_m_write
	wire    [4:0] dma_0_m_burstcount;                                               // dma_0:m_burstcount -> mm_interconnect_3:dma_0_m_burstcount
	wire  [511:0] mm_interconnect_3_clock_cross_dma_to_pcie_s0_readdata;            // clock_cross_dma_to_pcie:s0_readdata -> mm_interconnect_3:clock_cross_dma_to_pcie_s0_readdata
	wire          mm_interconnect_3_clock_cross_dma_to_pcie_s0_waitrequest;         // clock_cross_dma_to_pcie:s0_waitrequest -> mm_interconnect_3:clock_cross_dma_to_pcie_s0_waitrequest
	wire          mm_interconnect_3_clock_cross_dma_to_pcie_s0_debugaccess;         // mm_interconnect_3:clock_cross_dma_to_pcie_s0_debugaccess -> clock_cross_dma_to_pcie:s0_debugaccess
	wire   [19:0] mm_interconnect_3_clock_cross_dma_to_pcie_s0_address;             // mm_interconnect_3:clock_cross_dma_to_pcie_s0_address -> clock_cross_dma_to_pcie:s0_address
	wire          mm_interconnect_3_clock_cross_dma_to_pcie_s0_read;                // mm_interconnect_3:clock_cross_dma_to_pcie_s0_read -> clock_cross_dma_to_pcie:s0_read
	wire   [63:0] mm_interconnect_3_clock_cross_dma_to_pcie_s0_byteenable;          // mm_interconnect_3:clock_cross_dma_to_pcie_s0_byteenable -> clock_cross_dma_to_pcie:s0_byteenable
	wire          mm_interconnect_3_clock_cross_dma_to_pcie_s0_readdatavalid;       // clock_cross_dma_to_pcie:s0_readdatavalid -> mm_interconnect_3:clock_cross_dma_to_pcie_s0_readdatavalid
	wire          mm_interconnect_3_clock_cross_dma_to_pcie_s0_write;               // mm_interconnect_3:clock_cross_dma_to_pcie_s0_write -> clock_cross_dma_to_pcie:s0_write
	wire  [511:0] mm_interconnect_3_clock_cross_dma_to_pcie_s0_writedata;           // mm_interconnect_3:clock_cross_dma_to_pcie_s0_writedata -> clock_cross_dma_to_pcie:s0_writedata
	wire    [4:0] mm_interconnect_3_clock_cross_dma_to_pcie_s0_burstcount;          // mm_interconnect_3:clock_cross_dma_to_pcie_s0_burstcount -> clock_cross_dma_to_pcie:s0_burstcount
	wire          mm_interconnect_3_acl_memory_bank_divider_0_s_beginbursttransfer; // mm_interconnect_3:acl_memory_bank_divider_0_s_beginbursttransfer -> acl_memory_bank_divider_0:s_beginbursttransfer
	wire  [511:0] mm_interconnect_3_acl_memory_bank_divider_0_s_readdata;           // acl_memory_bank_divider_0:s_readdata -> mm_interconnect_3:acl_memory_bank_divider_0_s_readdata
	wire          mm_interconnect_3_acl_memory_bank_divider_0_s_waitrequest;        // acl_memory_bank_divider_0:s_waitrequest -> mm_interconnect_3:acl_memory_bank_divider_0_s_waitrequest
	wire   [25:0] mm_interconnect_3_acl_memory_bank_divider_0_s_address;            // mm_interconnect_3:acl_memory_bank_divider_0_s_address -> acl_memory_bank_divider_0:s_address
	wire          mm_interconnect_3_acl_memory_bank_divider_0_s_read;               // mm_interconnect_3:acl_memory_bank_divider_0_s_read -> acl_memory_bank_divider_0:s_read
	wire   [63:0] mm_interconnect_3_acl_memory_bank_divider_0_s_byteenable;         // mm_interconnect_3:acl_memory_bank_divider_0_s_byteenable -> acl_memory_bank_divider_0:s_byteenable
	wire          mm_interconnect_3_acl_memory_bank_divider_0_s_readdatavalid;      // acl_memory_bank_divider_0:s_readdatavalid -> mm_interconnect_3:acl_memory_bank_divider_0_s_readdatavalid
	wire          mm_interconnect_3_acl_memory_bank_divider_0_s_write;              // mm_interconnect_3:acl_memory_bank_divider_0_s_write -> acl_memory_bank_divider_0:s_write
	wire  [511:0] mm_interconnect_3_acl_memory_bank_divider_0_s_writedata;          // mm_interconnect_3:acl_memory_bank_divider_0_s_writedata -> acl_memory_bank_divider_0:s_writedata
	wire    [4:0] mm_interconnect_3_acl_memory_bank_divider_0_s_burstcount;         // mm_interconnect_3:acl_memory_bank_divider_0_s_burstcount -> acl_memory_bank_divider_0:s_burstcount
	wire          clock_cross_kernel_mem_0_m0_waitrequest;                          // mm_interconnect_5:clock_cross_kernel_mem_0_m0_waitrequest -> clock_cross_kernel_mem_0:m0_waitrequest
	wire  [511:0] clock_cross_kernel_mem_0_m0_readdata;                             // mm_interconnect_5:clock_cross_kernel_mem_0_m0_readdata -> clock_cross_kernel_mem_0:m0_readdata
	wire          clock_cross_kernel_mem_0_m0_debugaccess;                          // clock_cross_kernel_mem_0:m0_debugaccess -> mm_interconnect_5:clock_cross_kernel_mem_0_m0_debugaccess
	wire   [30:0] clock_cross_kernel_mem_0_m0_address;                              // clock_cross_kernel_mem_0:m0_address -> mm_interconnect_5:clock_cross_kernel_mem_0_m0_address
	wire          clock_cross_kernel_mem_0_m0_read;                                 // clock_cross_kernel_mem_0:m0_read -> mm_interconnect_5:clock_cross_kernel_mem_0_m0_read
	wire   [63:0] clock_cross_kernel_mem_0_m0_byteenable;                           // clock_cross_kernel_mem_0:m0_byteenable -> mm_interconnect_5:clock_cross_kernel_mem_0_m0_byteenable
	wire          clock_cross_kernel_mem_0_m0_readdatavalid;                        // mm_interconnect_5:clock_cross_kernel_mem_0_m0_readdatavalid -> clock_cross_kernel_mem_0:m0_readdatavalid
	wire  [511:0] clock_cross_kernel_mem_0_m0_writedata;                            // clock_cross_kernel_mem_0:m0_writedata -> mm_interconnect_5:clock_cross_kernel_mem_0_m0_writedata
	wire          clock_cross_kernel_mem_0_m0_write;                                // clock_cross_kernel_mem_0:m0_write -> mm_interconnect_5:clock_cross_kernel_mem_0_m0_write
	wire    [4:0] clock_cross_kernel_mem_0_m0_burstcount;                           // clock_cross_kernel_mem_0:m0_burstcount -> mm_interconnect_5:clock_cross_kernel_mem_0_m0_burstcount
	wire          mm_interconnect_5_em_pc_0_avl_in_beginbursttransfer;              // mm_interconnect_5:em_pc_0_avl_in_beginbursttransfer -> em_pc_0:avl_in_beginbursttransfer
	wire  [511:0] mm_interconnect_5_em_pc_0_avl_in_readdata;                        // em_pc_0:avl_in_readdata -> mm_interconnect_5:em_pc_0_avl_in_readdata
	wire          mm_interconnect_5_em_pc_0_avl_in_waitrequest;                     // em_pc_0:avl_in_waitrequest -> mm_interconnect_5:em_pc_0_avl_in_waitrequest
	wire   [24:0] mm_interconnect_5_em_pc_0_avl_in_address;                         // mm_interconnect_5:em_pc_0_avl_in_address -> em_pc_0:avl_in_address
	wire          mm_interconnect_5_em_pc_0_avl_in_read;                            // mm_interconnect_5:em_pc_0_avl_in_read -> em_pc_0:avl_in_read
	wire   [63:0] mm_interconnect_5_em_pc_0_avl_in_byteenable;                      // mm_interconnect_5:em_pc_0_avl_in_byteenable -> em_pc_0:avl_in_byteenable
	wire          mm_interconnect_5_em_pc_0_avl_in_readdatavalid;                   // em_pc_0:avl_in_readdatavalid -> mm_interconnect_5:em_pc_0_avl_in_readdatavalid
	wire          mm_interconnect_5_em_pc_0_avl_in_write;                           // mm_interconnect_5:em_pc_0_avl_in_write -> em_pc_0:avl_in_write
	wire  [511:0] mm_interconnect_5_em_pc_0_avl_in_writedata;                       // mm_interconnect_5:em_pc_0_avl_in_writedata -> em_pc_0:avl_in_writedata
	wire    [0:0] mm_interconnect_5_em_pc_0_avl_in_burstcount;                      // mm_interconnect_5:em_pc_0_avl_in_burstcount -> em_pc_0:avl_in_burstcount
	wire          em_pc_0_avl_out_beginbursttransfer;                               // em_pc_0:avl_out_beginbursttransfer -> mm_interconnect_6:em_pc_0_avl_out_beginbursttransfer
	wire          em_pc_0_avl_out_waitrequest;                                      // mm_interconnect_6:em_pc_0_avl_out_waitrequest -> em_pc_0:avl_out_waitrequest
	wire  [511:0] em_pc_0_avl_out_readdata;                                         // mm_interconnect_6:em_pc_0_avl_out_readdata -> em_pc_0:avl_out_readdata
	wire   [30:0] em_pc_0_avl_out_address;                                          // em_pc_0:avl_out_address -> mm_interconnect_6:em_pc_0_avl_out_address
	wire   [63:0] em_pc_0_avl_out_byteenable;                                       // em_pc_0:avl_out_byteenable -> mm_interconnect_6:em_pc_0_avl_out_byteenable
	wire          em_pc_0_avl_out_read;                                             // em_pc_0:avl_out_read -> mm_interconnect_6:em_pc_0_avl_out_read
	wire          em_pc_0_avl_out_readdatavalid;                                    // mm_interconnect_6:em_pc_0_avl_out_readdatavalid -> em_pc_0:avl_out_readdatavalid
	wire          em_pc_0_avl_out_write;                                            // em_pc_0:avl_out_write -> mm_interconnect_6:em_pc_0_avl_out_write
	wire  [511:0] em_pc_0_avl_out_writedata;                                        // em_pc_0:avl_out_writedata -> mm_interconnect_6:em_pc_0_avl_out_writedata
	wire          em_pc_0_avl_out_burstcount;                                       // em_pc_0:avl_out_burstcount -> mm_interconnect_6:em_pc_0_avl_out_burstcount
	wire          acl_memory_bank_divider_0_bank1_waitrequest;                      // mm_interconnect_6:acl_memory_bank_divider_0_bank1_waitrequest -> acl_memory_bank_divider_0:bank1_waitrequest
	wire  [511:0] acl_memory_bank_divider_0_bank1_readdata;                         // mm_interconnect_6:acl_memory_bank_divider_0_bank1_readdata -> acl_memory_bank_divider_0:bank1_readdata
	wire   [30:0] acl_memory_bank_divider_0_bank1_address;                          // acl_memory_bank_divider_0:bank1_address -> mm_interconnect_6:acl_memory_bank_divider_0_bank1_address
	wire          acl_memory_bank_divider_0_bank1_read;                             // acl_memory_bank_divider_0:bank1_read -> mm_interconnect_6:acl_memory_bank_divider_0_bank1_read
	wire   [63:0] acl_memory_bank_divider_0_bank1_byteenable;                       // acl_memory_bank_divider_0:bank1_byteenable -> mm_interconnect_6:acl_memory_bank_divider_0_bank1_byteenable
	wire          acl_memory_bank_divider_0_bank1_readdatavalid;                    // mm_interconnect_6:acl_memory_bank_divider_0_bank1_readdatavalid -> acl_memory_bank_divider_0:bank1_readdatavalid
	wire  [511:0] acl_memory_bank_divider_0_bank1_writedata;                        // acl_memory_bank_divider_0:bank1_writedata -> mm_interconnect_6:acl_memory_bank_divider_0_bank1_writedata
	wire          acl_memory_bank_divider_0_bank1_write;                            // acl_memory_bank_divider_0:bank1_write -> mm_interconnect_6:acl_memory_bank_divider_0_bank1_write
	wire    [4:0] acl_memory_bank_divider_0_bank1_burstcount;                       // acl_memory_bank_divider_0:bank1_burstcount -> mm_interconnect_6:acl_memory_bank_divider_0_bank1_burstcount
	wire  [511:0] mm_interconnect_6_pipe_stage_ddr3a_iface_s0_readdata;             // pipe_stage_ddr3a_iface:s0_readdata -> mm_interconnect_6:pipe_stage_ddr3a_iface_s0_readdata
	wire          mm_interconnect_6_pipe_stage_ddr3a_iface_s0_waitrequest;          // pipe_stage_ddr3a_iface:s0_waitrequest -> mm_interconnect_6:pipe_stage_ddr3a_iface_s0_waitrequest
	wire          mm_interconnect_6_pipe_stage_ddr3a_iface_s0_debugaccess;          // mm_interconnect_6:pipe_stage_ddr3a_iface_s0_debugaccess -> pipe_stage_ddr3a_iface:s0_debugaccess
	wire   [30:0] mm_interconnect_6_pipe_stage_ddr3a_iface_s0_address;              // mm_interconnect_6:pipe_stage_ddr3a_iface_s0_address -> pipe_stage_ddr3a_iface:s0_address
	wire          mm_interconnect_6_pipe_stage_ddr3a_iface_s0_read;                 // mm_interconnect_6:pipe_stage_ddr3a_iface_s0_read -> pipe_stage_ddr3a_iface:s0_read
	wire   [63:0] mm_interconnect_6_pipe_stage_ddr3a_iface_s0_byteenable;           // mm_interconnect_6:pipe_stage_ddr3a_iface_s0_byteenable -> pipe_stage_ddr3a_iface:s0_byteenable
	wire          mm_interconnect_6_pipe_stage_ddr3a_iface_s0_readdatavalid;        // pipe_stage_ddr3a_iface:s0_readdatavalid -> mm_interconnect_6:pipe_stage_ddr3a_iface_s0_readdatavalid
	wire          mm_interconnect_6_pipe_stage_ddr3a_iface_s0_write;                // mm_interconnect_6:pipe_stage_ddr3a_iface_s0_write -> pipe_stage_ddr3a_iface:s0_write
	wire  [511:0] mm_interconnect_6_pipe_stage_ddr3a_iface_s0_writedata;            // mm_interconnect_6:pipe_stage_ddr3a_iface_s0_writedata -> pipe_stage_ddr3a_iface:s0_writedata
	wire    [4:0] mm_interconnect_6_pipe_stage_ddr3a_iface_s0_burstcount;           // mm_interconnect_6:pipe_stage_ddr3a_iface_s0_burstcount -> pipe_stage_ddr3a_iface:s0_burstcount
	wire          clock_cross_kernel_mem_1_m0_waitrequest;                          // mm_interconnect_7:clock_cross_kernel_mem_1_m0_waitrequest -> clock_cross_kernel_mem_1:m0_waitrequest
	wire  [511:0] clock_cross_kernel_mem_1_m0_readdata;                             // mm_interconnect_7:clock_cross_kernel_mem_1_m0_readdata -> clock_cross_kernel_mem_1:m0_readdata
	wire          clock_cross_kernel_mem_1_m0_debugaccess;                          // clock_cross_kernel_mem_1:m0_debugaccess -> mm_interconnect_7:clock_cross_kernel_mem_1_m0_debugaccess
	wire   [30:0] clock_cross_kernel_mem_1_m0_address;                              // clock_cross_kernel_mem_1:m0_address -> mm_interconnect_7:clock_cross_kernel_mem_1_m0_address
	wire          clock_cross_kernel_mem_1_m0_read;                                 // clock_cross_kernel_mem_1:m0_read -> mm_interconnect_7:clock_cross_kernel_mem_1_m0_read
	wire   [63:0] clock_cross_kernel_mem_1_m0_byteenable;                           // clock_cross_kernel_mem_1:m0_byteenable -> mm_interconnect_7:clock_cross_kernel_mem_1_m0_byteenable
	wire          clock_cross_kernel_mem_1_m0_readdatavalid;                        // mm_interconnect_7:clock_cross_kernel_mem_1_m0_readdatavalid -> clock_cross_kernel_mem_1:m0_readdatavalid
	wire  [511:0] clock_cross_kernel_mem_1_m0_writedata;                            // clock_cross_kernel_mem_1:m0_writedata -> mm_interconnect_7:clock_cross_kernel_mem_1_m0_writedata
	wire          clock_cross_kernel_mem_1_m0_write;                                // clock_cross_kernel_mem_1:m0_write -> mm_interconnect_7:clock_cross_kernel_mem_1_m0_write
	wire    [4:0] clock_cross_kernel_mem_1_m0_burstcount;                           // clock_cross_kernel_mem_1:m0_burstcount -> mm_interconnect_7:clock_cross_kernel_mem_1_m0_burstcount
	wire          mm_interconnect_7_em_pc_1_avl_in_beginbursttransfer;              // mm_interconnect_7:em_pc_1_avl_in_beginbursttransfer -> em_pc_1:avl_in_beginbursttransfer
	wire  [511:0] mm_interconnect_7_em_pc_1_avl_in_readdata;                        // em_pc_1:avl_in_readdata -> mm_interconnect_7:em_pc_1_avl_in_readdata
	wire          mm_interconnect_7_em_pc_1_avl_in_waitrequest;                     // em_pc_1:avl_in_waitrequest -> mm_interconnect_7:em_pc_1_avl_in_waitrequest
	wire   [24:0] mm_interconnect_7_em_pc_1_avl_in_address;                         // mm_interconnect_7:em_pc_1_avl_in_address -> em_pc_1:avl_in_address
	wire          mm_interconnect_7_em_pc_1_avl_in_read;                            // mm_interconnect_7:em_pc_1_avl_in_read -> em_pc_1:avl_in_read
	wire   [63:0] mm_interconnect_7_em_pc_1_avl_in_byteenable;                      // mm_interconnect_7:em_pc_1_avl_in_byteenable -> em_pc_1:avl_in_byteenable
	wire          mm_interconnect_7_em_pc_1_avl_in_readdatavalid;                   // em_pc_1:avl_in_readdatavalid -> mm_interconnect_7:em_pc_1_avl_in_readdatavalid
	wire          mm_interconnect_7_em_pc_1_avl_in_write;                           // mm_interconnect_7:em_pc_1_avl_in_write -> em_pc_1:avl_in_write
	wire  [511:0] mm_interconnect_7_em_pc_1_avl_in_writedata;                       // mm_interconnect_7:em_pc_1_avl_in_writedata -> em_pc_1:avl_in_writedata
	wire    [0:0] mm_interconnect_7_em_pc_1_avl_in_burstcount;                      // mm_interconnect_7:em_pc_1_avl_in_burstcount -> em_pc_1:avl_in_burstcount
	wire          pcie_rxm_bar0_waitrequest;                                        // mm_interconnect_8:pcie_Rxm_BAR0_waitrequest -> pcie:RxmWaitRequest_0_i
	wire  [127:0] pcie_rxm_bar0_readdata;                                           // mm_interconnect_8:pcie_Rxm_BAR0_readdata -> pcie:RxmReadData_0_i
	wire   [31:0] pcie_rxm_bar0_address;                                            // pcie:RxmAddress_0_o -> mm_interconnect_8:pcie_Rxm_BAR0_address
	wire          pcie_rxm_bar0_read;                                               // pcie:RxmRead_0_o -> mm_interconnect_8:pcie_Rxm_BAR0_read
	wire   [15:0] pcie_rxm_bar0_byteenable;                                         // pcie:RxmByteEnable_0_o -> mm_interconnect_8:pcie_Rxm_BAR0_byteenable
	wire          pcie_rxm_bar0_readdatavalid;                                      // mm_interconnect_8:pcie_Rxm_BAR0_readdatavalid -> pcie:RxmReadDataValid_0_i
	wire          pcie_rxm_bar0_write;                                              // pcie:RxmWrite_0_o -> mm_interconnect_8:pcie_Rxm_BAR0_write
	wire  [127:0] pcie_rxm_bar0_writedata;                                          // pcie:RxmWriteData_0_o -> mm_interconnect_8:pcie_Rxm_BAR0_writedata
	wire    [5:0] pcie_rxm_bar0_burstcount;                                         // pcie:RxmBurstCount_0_o -> mm_interconnect_8:pcie_Rxm_BAR0_burstcount
	wire   [31:0] mm_interconnect_8_pipe_stage_host_ctrl_s0_readdata;               // pipe_stage_host_ctrl:s0_readdata -> mm_interconnect_8:pipe_stage_host_ctrl_s0_readdata
	wire          mm_interconnect_8_pipe_stage_host_ctrl_s0_waitrequest;            // pipe_stage_host_ctrl:s0_waitrequest -> mm_interconnect_8:pipe_stage_host_ctrl_s0_waitrequest
	wire          mm_interconnect_8_pipe_stage_host_ctrl_s0_debugaccess;            // mm_interconnect_8:pipe_stage_host_ctrl_s0_debugaccess -> pipe_stage_host_ctrl:s0_debugaccess
	wire   [17:0] mm_interconnect_8_pipe_stage_host_ctrl_s0_address;                // mm_interconnect_8:pipe_stage_host_ctrl_s0_address -> pipe_stage_host_ctrl:s0_address
	wire          mm_interconnect_8_pipe_stage_host_ctrl_s0_read;                   // mm_interconnect_8:pipe_stage_host_ctrl_s0_read -> pipe_stage_host_ctrl:s0_read
	wire    [3:0] mm_interconnect_8_pipe_stage_host_ctrl_s0_byteenable;             // mm_interconnect_8:pipe_stage_host_ctrl_s0_byteenable -> pipe_stage_host_ctrl:s0_byteenable
	wire          mm_interconnect_8_pipe_stage_host_ctrl_s0_readdatavalid;          // pipe_stage_host_ctrl:s0_readdatavalid -> mm_interconnect_8:pipe_stage_host_ctrl_s0_readdatavalid
	wire          mm_interconnect_8_pipe_stage_host_ctrl_s0_write;                  // mm_interconnect_8:pipe_stage_host_ctrl_s0_write -> pipe_stage_host_ctrl:s0_write
	wire   [31:0] mm_interconnect_8_pipe_stage_host_ctrl_s0_writedata;              // mm_interconnect_8:pipe_stage_host_ctrl_s0_writedata -> pipe_stage_host_ctrl:s0_writedata
	wire    [0:0] mm_interconnect_8_pipe_stage_host_ctrl_s0_burstcount;             // mm_interconnect_8:pipe_stage_host_ctrl_s0_burstcount -> pipe_stage_host_ctrl:s0_burstcount
	wire          clock_cross_dma_to_pcie_m0_waitrequest;                           // mm_interconnect_9:clock_cross_dma_to_pcie_m0_waitrequest -> clock_cross_dma_to_pcie:m0_waitrequest
	wire  [511:0] clock_cross_dma_to_pcie_m0_readdata;                              // mm_interconnect_9:clock_cross_dma_to_pcie_m0_readdata -> clock_cross_dma_to_pcie:m0_readdata
	wire          clock_cross_dma_to_pcie_m0_debugaccess;                           // clock_cross_dma_to_pcie:m0_debugaccess -> mm_interconnect_9:clock_cross_dma_to_pcie_m0_debugaccess
	wire   [19:0] clock_cross_dma_to_pcie_m0_address;                               // clock_cross_dma_to_pcie:m0_address -> mm_interconnect_9:clock_cross_dma_to_pcie_m0_address
	wire          clock_cross_dma_to_pcie_m0_read;                                  // clock_cross_dma_to_pcie:m0_read -> mm_interconnect_9:clock_cross_dma_to_pcie_m0_read
	wire   [63:0] clock_cross_dma_to_pcie_m0_byteenable;                            // clock_cross_dma_to_pcie:m0_byteenable -> mm_interconnect_9:clock_cross_dma_to_pcie_m0_byteenable
	wire          clock_cross_dma_to_pcie_m0_readdatavalid;                         // mm_interconnect_9:clock_cross_dma_to_pcie_m0_readdatavalid -> clock_cross_dma_to_pcie:m0_readdatavalid
	wire  [511:0] clock_cross_dma_to_pcie_m0_writedata;                             // clock_cross_dma_to_pcie:m0_writedata -> mm_interconnect_9:clock_cross_dma_to_pcie_m0_writedata
	wire          clock_cross_dma_to_pcie_m0_write;                                 // clock_cross_dma_to_pcie:m0_write -> mm_interconnect_9:clock_cross_dma_to_pcie_m0_write
	wire    [4:0] clock_cross_dma_to_pcie_m0_burstcount;                            // clock_cross_dma_to_pcie:m0_burstcount -> mm_interconnect_9:clock_cross_dma_to_pcie_m0_burstcount
	wire          mm_interconnect_9_pcie_txs_chipselect;                            // mm_interconnect_9:pcie_Txs_chipselect -> pcie:TxsChipSelect_i
	wire  [127:0] mm_interconnect_9_pcie_txs_readdata;                              // pcie:TxsReadData_o -> mm_interconnect_9:pcie_Txs_readdata
	wire          mm_interconnect_9_pcie_txs_waitrequest;                           // pcie:TxsWaitRequest_o -> mm_interconnect_9:pcie_Txs_waitrequest
	wire   [19:0] mm_interconnect_9_pcie_txs_address;                               // mm_interconnect_9:pcie_Txs_address -> pcie:TxsAddress_i
	wire          mm_interconnect_9_pcie_txs_read;                                  // mm_interconnect_9:pcie_Txs_read -> pcie:TxsRead_i
	wire   [15:0] mm_interconnect_9_pcie_txs_byteenable;                            // mm_interconnect_9:pcie_Txs_byteenable -> pcie:TxsByteEnable_i
	wire          mm_interconnect_9_pcie_txs_readdatavalid;                         // pcie:TxsReadDataValid_o -> mm_interconnect_9:pcie_Txs_readdatavalid
	wire          mm_interconnect_9_pcie_txs_write;                                 // mm_interconnect_9:pcie_Txs_write -> pcie:TxsWrite_i
	wire  [127:0] mm_interconnect_9_pcie_txs_writedata;                             // mm_interconnect_9:pcie_Txs_writedata -> pcie:TxsWriteData_i
	wire    [5:0] mm_interconnect_9_pcie_txs_burstcount;                            // mm_interconnect_9:pcie_Txs_burstcount -> pcie:TxsBurstCount_i
	wire          em_pc_1_avl_out_beginbursttransfer;                               // em_pc_1:avl_out_beginbursttransfer -> mm_interconnect_10:em_pc_1_avl_out_beginbursttransfer
	wire          em_pc_1_avl_out_waitrequest;                                      // mm_interconnect_10:em_pc_1_avl_out_waitrequest -> em_pc_1:avl_out_waitrequest
	wire  [511:0] em_pc_1_avl_out_readdata;                                         // mm_interconnect_10:em_pc_1_avl_out_readdata -> em_pc_1:avl_out_readdata
	wire   [30:0] em_pc_1_avl_out_address;                                          // em_pc_1:avl_out_address -> mm_interconnect_10:em_pc_1_avl_out_address
	wire   [63:0] em_pc_1_avl_out_byteenable;                                       // em_pc_1:avl_out_byteenable -> mm_interconnect_10:em_pc_1_avl_out_byteenable
	wire          em_pc_1_avl_out_read;                                             // em_pc_1:avl_out_read -> mm_interconnect_10:em_pc_1_avl_out_read
	wire          em_pc_1_avl_out_readdatavalid;                                    // mm_interconnect_10:em_pc_1_avl_out_readdatavalid -> em_pc_1:avl_out_readdatavalid
	wire          em_pc_1_avl_out_write;                                            // em_pc_1:avl_out_write -> mm_interconnect_10:em_pc_1_avl_out_write
	wire  [511:0] em_pc_1_avl_out_writedata;                                        // em_pc_1:avl_out_writedata -> mm_interconnect_10:em_pc_1_avl_out_writedata
	wire          em_pc_1_avl_out_burstcount;                                       // em_pc_1:avl_out_burstcount -> mm_interconnect_10:em_pc_1_avl_out_burstcount
	wire          clock_cross_dma_to_ddr3b_m0_waitrequest;                          // mm_interconnect_10:clock_cross_dma_to_ddr3b_m0_waitrequest -> clock_cross_dma_to_ddr3b:m0_waitrequest
	wire  [511:0] clock_cross_dma_to_ddr3b_m0_readdata;                             // mm_interconnect_10:clock_cross_dma_to_ddr3b_m0_readdata -> clock_cross_dma_to_ddr3b:m0_readdata
	wire          clock_cross_dma_to_ddr3b_m0_debugaccess;                          // clock_cross_dma_to_ddr3b:m0_debugaccess -> mm_interconnect_10:clock_cross_dma_to_ddr3b_m0_debugaccess
	wire   [30:0] clock_cross_dma_to_ddr3b_m0_address;                              // clock_cross_dma_to_ddr3b:m0_address -> mm_interconnect_10:clock_cross_dma_to_ddr3b_m0_address
	wire          clock_cross_dma_to_ddr3b_m0_read;                                 // clock_cross_dma_to_ddr3b:m0_read -> mm_interconnect_10:clock_cross_dma_to_ddr3b_m0_read
	wire   [63:0] clock_cross_dma_to_ddr3b_m0_byteenable;                           // clock_cross_dma_to_ddr3b:m0_byteenable -> mm_interconnect_10:clock_cross_dma_to_ddr3b_m0_byteenable
	wire          clock_cross_dma_to_ddr3b_m0_readdatavalid;                        // mm_interconnect_10:clock_cross_dma_to_ddr3b_m0_readdatavalid -> clock_cross_dma_to_ddr3b:m0_readdatavalid
	wire  [511:0] clock_cross_dma_to_ddr3b_m0_writedata;                            // clock_cross_dma_to_ddr3b:m0_writedata -> mm_interconnect_10:clock_cross_dma_to_ddr3b_m0_writedata
	wire          clock_cross_dma_to_ddr3b_m0_write;                                // clock_cross_dma_to_ddr3b:m0_write -> mm_interconnect_10:clock_cross_dma_to_ddr3b_m0_write
	wire    [4:0] clock_cross_dma_to_ddr3b_m0_burstcount;                           // clock_cross_dma_to_ddr3b:m0_burstcount -> mm_interconnect_10:clock_cross_dma_to_ddr3b_m0_burstcount
	wire  [511:0] mm_interconnect_10_pipe_stage_ddr3b_iface_s0_readdata;            // pipe_stage_ddr3b_iface:s0_readdata -> mm_interconnect_10:pipe_stage_ddr3b_iface_s0_readdata
	wire          mm_interconnect_10_pipe_stage_ddr3b_iface_s0_waitrequest;         // pipe_stage_ddr3b_iface:s0_waitrequest -> mm_interconnect_10:pipe_stage_ddr3b_iface_s0_waitrequest
	wire          mm_interconnect_10_pipe_stage_ddr3b_iface_s0_debugaccess;         // mm_interconnect_10:pipe_stage_ddr3b_iface_s0_debugaccess -> pipe_stage_ddr3b_iface:s0_debugaccess
	wire   [30:0] mm_interconnect_10_pipe_stage_ddr3b_iface_s0_address;             // mm_interconnect_10:pipe_stage_ddr3b_iface_s0_address -> pipe_stage_ddr3b_iface:s0_address
	wire          mm_interconnect_10_pipe_stage_ddr3b_iface_s0_read;                // mm_interconnect_10:pipe_stage_ddr3b_iface_s0_read -> pipe_stage_ddr3b_iface:s0_read
	wire   [63:0] mm_interconnect_10_pipe_stage_ddr3b_iface_s0_byteenable;          // mm_interconnect_10:pipe_stage_ddr3b_iface_s0_byteenable -> pipe_stage_ddr3b_iface:s0_byteenable
	wire          mm_interconnect_10_pipe_stage_ddr3b_iface_s0_readdatavalid;       // pipe_stage_ddr3b_iface:s0_readdatavalid -> mm_interconnect_10:pipe_stage_ddr3b_iface_s0_readdatavalid
	wire          mm_interconnect_10_pipe_stage_ddr3b_iface_s0_write;               // mm_interconnect_10:pipe_stage_ddr3b_iface_s0_write -> pipe_stage_ddr3b_iface:s0_write
	wire  [511:0] mm_interconnect_10_pipe_stage_ddr3b_iface_s0_writedata;           // mm_interconnect_10:pipe_stage_ddr3b_iface_s0_writedata -> pipe_stage_ddr3b_iface:s0_writedata
	wire    [4:0] mm_interconnect_10_pipe_stage_ddr3b_iface_s0_burstcount;          // mm_interconnect_10:pipe_stage_ddr3b_iface_s0_burstcount -> pipe_stage_ddr3b_iface:s0_burstcount
	wire          acl_memory_bank_divider_0_bank2_waitrequest;                      // mm_interconnect_12:acl_memory_bank_divider_0_bank2_waitrequest -> acl_memory_bank_divider_0:bank2_waitrequest
	wire  [511:0] acl_memory_bank_divider_0_bank2_readdata;                         // mm_interconnect_12:acl_memory_bank_divider_0_bank2_readdata -> acl_memory_bank_divider_0:bank2_readdata
	wire   [30:0] acl_memory_bank_divider_0_bank2_address;                          // acl_memory_bank_divider_0:bank2_address -> mm_interconnect_12:acl_memory_bank_divider_0_bank2_address
	wire          acl_memory_bank_divider_0_bank2_read;                             // acl_memory_bank_divider_0:bank2_read -> mm_interconnect_12:acl_memory_bank_divider_0_bank2_read
	wire   [63:0] acl_memory_bank_divider_0_bank2_byteenable;                       // acl_memory_bank_divider_0:bank2_byteenable -> mm_interconnect_12:acl_memory_bank_divider_0_bank2_byteenable
	wire          acl_memory_bank_divider_0_bank2_readdatavalid;                    // mm_interconnect_12:acl_memory_bank_divider_0_bank2_readdatavalid -> acl_memory_bank_divider_0:bank2_readdatavalid
	wire  [511:0] acl_memory_bank_divider_0_bank2_writedata;                        // acl_memory_bank_divider_0:bank2_writedata -> mm_interconnect_12:acl_memory_bank_divider_0_bank2_writedata
	wire          acl_memory_bank_divider_0_bank2_write;                            // acl_memory_bank_divider_0:bank2_write -> mm_interconnect_12:acl_memory_bank_divider_0_bank2_write
	wire    [4:0] acl_memory_bank_divider_0_bank2_burstcount;                       // acl_memory_bank_divider_0:bank2_burstcount -> mm_interconnect_12:acl_memory_bank_divider_0_bank2_burstcount
	wire  [511:0] mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_readdata;          // clock_cross_dma_to_ddr3b:s0_readdata -> mm_interconnect_12:clock_cross_dma_to_ddr3b_s0_readdata
	wire          mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_waitrequest;       // clock_cross_dma_to_ddr3b:s0_waitrequest -> mm_interconnect_12:clock_cross_dma_to_ddr3b_s0_waitrequest
	wire          mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_debugaccess;       // mm_interconnect_12:clock_cross_dma_to_ddr3b_s0_debugaccess -> clock_cross_dma_to_ddr3b:s0_debugaccess
	wire   [30:0] mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_address;           // mm_interconnect_12:clock_cross_dma_to_ddr3b_s0_address -> clock_cross_dma_to_ddr3b:s0_address
	wire          mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_read;              // mm_interconnect_12:clock_cross_dma_to_ddr3b_s0_read -> clock_cross_dma_to_ddr3b:s0_read
	wire   [63:0] mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_byteenable;        // mm_interconnect_12:clock_cross_dma_to_ddr3b_s0_byteenable -> clock_cross_dma_to_ddr3b:s0_byteenable
	wire          mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_readdatavalid;     // clock_cross_dma_to_ddr3b:s0_readdatavalid -> mm_interconnect_12:clock_cross_dma_to_ddr3b_s0_readdatavalid
	wire          mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_write;             // mm_interconnect_12:clock_cross_dma_to_ddr3b_s0_write -> clock_cross_dma_to_ddr3b:s0_write
	wire  [511:0] mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_writedata;         // mm_interconnect_12:clock_cross_dma_to_ddr3b_s0_writedata -> clock_cross_dma_to_ddr3b:s0_writedata
	wire    [4:0] mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_burstcount;        // mm_interconnect_12:clock_cross_dma_to_ddr3b_s0_burstcount -> clock_cross_dma_to_ddr3b:s0_burstcount
	wire   [15:0] pcie_rxmirq_irq;                                                  // irq_mapper:sender_irq -> pcie:RxmIrq_i
	wire          irq_mapper_receiver0_irq;                                         // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                    // kernel_interface:kernel_irq_to_host_irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver1_irq;                                         // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                // dma_0:dma_irq_irq -> irq_synchronizer_001:receiver_irq
	wire          rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [clock_cross_dma_to_pcie:s0_reset, mm_interconnect_0:ddr3a_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:ddr3a_soft_reset_reset_bridge_in_reset_reset, mm_interconnect_3:clock_cross_dma_to_pcie_s0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                               // rst_controller_001:reset_out -> [mm_interconnect_2:temperature_0_clk_reset_reset_bridge_in_reset_reset, temperature_0:resetn]
	wire          rst_controller_002_reset_out_reset;                               // rst_controller_002:reset_out -> [acl_memory_bank_divider_0:reset_reset_n, dma_0:reset_reset_n, irq_synchronizer_001:receiver_reset, mm_interconnect_12:acl_memory_bank_divider_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:dma_0_reset_reset_bridge_in_reset_reset, mm_interconnect_3:dma_0_reset_reset_bridge_in_reset_reset, mm_interconnect_6:acl_memory_bank_divider_0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_003_reset_out_reset;                               // rst_controller_003:reset_out -> [clock_cross_kernel_mem_0:m0_reset, mm_interconnect_5:clock_cross_kernel_mem_0_m0_reset_reset_bridge_in_reset_reset]
	wire          kernel_interface_sw_reset_export_reset;                           // kernel_interface:sw_reset_export_reset_n -> [rst_controller_003:reset_in0, rst_controller_004:reset_in0]
	wire          rst_controller_004_reset_out_reset;                               // rst_controller_004:reset_out -> [clock_cross_kernel_mem_1:m0_reset, mm_interconnect_7:clock_cross_kernel_mem_1_m0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_005_reset_out_reset;                               // rst_controller_005:reset_out -> por_reset_counter:resetn
	wire          rst_controller_006_reset_out_reset;                               // rst_controller_006:reset_out -> [mm_interconnect_2:uniphy_status_0_clk_reset_reset_bridge_in_reset_reset, uniphy_status_0:resetn, version_id_0:resetn]
	wire          rst_controller_007_reset_out_reset;                               // rst_controller_007:reset_out -> [mm_interconnect_1:ddr3b_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ddr3b_soft_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_008_reset_out_reset;                               // rst_controller_008:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_2:pcie_Cra_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_8:pcie_Rxm_BAR0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_9:pcie_Txs_translator_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_009_reset_out_reset;                               // rst_controller_009:reset_out -> irq_synchronizer:receiver_reset

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (512),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (31),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pipe_stage_ddr3b_dimm (
		.clk              (ddr3b_afi_clk_clk),                       //   clk.clk
		.reset            (reset_controller_ddr3b_reset_out_reset),  // reset.reset
		.s0_waitrequest   (pipe_stage_ddr3b_iface_m0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (pipe_stage_ddr3b_iface_m0_readdata),      //      .readdata
		.s0_readdatavalid (pipe_stage_ddr3b_iface_m0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (pipe_stage_ddr3b_iface_m0_burstcount),    //      .burstcount
		.s0_writedata     (pipe_stage_ddr3b_iface_m0_writedata),     //      .writedata
		.s0_address       (pipe_stage_ddr3b_iface_m0_address),       //      .address
		.s0_write         (pipe_stage_ddr3b_iface_m0_write),         //      .write
		.s0_read          (pipe_stage_ddr3b_iface_m0_read),          //      .read
		.s0_byteenable    (pipe_stage_ddr3b_iface_m0_byteenable),    //      .byteenable
		.s0_debugaccess   (pipe_stage_ddr3b_iface_m0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pipe_stage_ddr3b_dimm_m0_waitrequest),    //    m0.waitrequest
		.m0_readdata      (pipe_stage_ddr3b_dimm_m0_readdata),       //      .readdata
		.m0_readdatavalid (pipe_stage_ddr3b_dimm_m0_readdatavalid),  //      .readdatavalid
		.m0_burstcount    (pipe_stage_ddr3b_dimm_m0_burstcount),     //      .burstcount
		.m0_writedata     (pipe_stage_ddr3b_dimm_m0_writedata),      //      .writedata
		.m0_address       (pipe_stage_ddr3b_dimm_m0_address),        //      .address
		.m0_write         (pipe_stage_ddr3b_dimm_m0_write),          //      .write
		.m0_read          (pipe_stage_ddr3b_dimm_m0_read),           //      .read
		.m0_byteenable    (pipe_stage_ddr3b_dimm_m0_byteenable),     //      .byteenable
		.m0_debugaccess   (pipe_stage_ddr3b_dimm_m0_debugaccess),    //      .debugaccess
		.s0_response      (),                                        // (terminated)
		.m0_response      (2'b00)                                    // (terminated)
	);

	altpcie_sv_hip_avmm_hwtcl #(
		.lane_mask_hwtcl                          ("x8"),
		.gen123_lane_rate_mode_hwtcl              ("Gen2 (5.0 Gbps)"),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("2.1"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.in_cvp_mode_hwtcl                        (1),
		.enable_tl_only_sim_hwtcl                 (0),
		.use_atx_pll_hwtcl                        (0),
		.enable_power_on_rst_pulse_hwtcl          (0),
		.enable_pcisigtest_hwtcl                  (0),
		.bar0_size_mask_hwtcl                     (18),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Enabled"),
		.bar0_prefetchable_hwtcl                  ("Enabled"),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_size_mask_hwtcl                     (0),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Disabled"),
		.bar2_prefetchable_hwtcl                  ("Disabled"),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_size_mask_hwtcl                     (0),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Disabled"),
		.bar4_prefetchable_hwtcl                  ("Disabled"),
		.bar5_size_mask_hwtcl                     (0),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.vendor_id_hwtcl                          (4466),
		.device_id_hwtcl                          (43776),
		.revision_id_hwtcl                        (1),
		.class_code_hwtcl                         (16711680),
		.subsystem_vendor_id_hwtcl                (4466),
		.subsystem_device_id_hwtcl                (4),
		.max_payload_size_hwtcl                   (256),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("ABCD"),
		.enable_completion_timeout_disable_hwtcl  (1),
		.use_aer_hwtcl                            (0),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("4"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.vsec_id_hwtcl                            (40960),
		.vsec_rev_hwtcl                           (0),
		.user_id_hwtcl                            (0),
		.avmm_width_hwtcl                         (128),
		.AVALON_ADDR_WIDTH                        (32),
		.avmm_burst_width_hwtcl                   (6),
		.CB_PCIE_MODE                             (0),
		.CB_PCIE_RX_LITE                          (0),
		.CB_RXM_DATA_WIDTH                        (128),
		.CG_AVALON_S_ADDR_WIDTH                   (20),
		.CG_IMPL_CRA_AV_SLAVE_PORT                (1),
		.CG_ENABLE_ADVANCED_INTERRUPT             (0),
		.CG_ENABLE_A2P_INTERRUPT                  (0),
		.CB_A2P_ADDR_MAP_IS_FIXED                 (0),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES              (256),
		.BYPASSS_A2P_TRANSLATION                  (0),
		.a2p_pass_thru_bits                       (12),
		.ast_width_hwtcl                          ("Avalon-ST 128-bit"),
		.use_ast_parity                           (0),
		.millisecond_cycle_count_hwtcl            (248500),
		.port_width_be_hwtcl                      (16),
		.port_width_data_hwtcl                    (128),
		.hip_reconfig_hwtcl                       (0),
		.expansion_base_address_register_hwtcl    (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.bypass_cdc_hwtcl                         ("false"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.device_number_hwtcl                      (0),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.maximum_current_hwtcl                    (0),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.disable_snoop_packet_hwtcl               ("false"),
		.enable_l1_aspm_hwtcl                     ("false"),
		.rx_ei_l0s_hwtcl                          (0),
		.enable_l0s_aspm_hwtcl                    ("false"),
		.aspm_config_management_hwtcl             ("true"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.extended_tag_reset_hwtcl                 ("false"),
		.no_command_completed_hwtcl               ("false"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.eie_before_nfts_count_hwtcl              (4),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("false"),
		.atomic_malformed_hwtcl                   ("true"),
		.flr_capability_hwtcl                     ("false"),
		.enable_adapter_half_rate_mode_hwtcl      ("false"),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("false"),
		.skp_os_gen3_count_hwtcl                  (0),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.retry_buffer_last_active_address_hwtcl   (2047),
		.reserved_debug_hwtcl                     (0),
		.bypass_clk_switch_hwtcl                  ("false"),
		.l2_async_logic_hwtcl                     ("disable"),
		.indicator_hwtcl                          (0),
		.diffclock_nfts_count_hwtcl               (128),
		.sameclock_nfts_count_hwtcl               (128),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.credit_buffer_allocation_aux_hwtcl       ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (195),
		.cpl_spc_data_hwtcl                       (781),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.cseb_cpl_status_during_cvp_hwtcl         ("completer_abort"),
		.core_clk_sel_hwtcl                       ("core_clk_250"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.g3_dis_rx_use_prst_hwtcl                 ("true"),
		.g3_dis_rx_use_prst_ep_hwtcl              ("true"),
		.deemphasis_enable_hwtcl                  ("false"),
		.reconfig_to_xcvr_width                   (700),
		.reconfig_from_xcvr_width                 (460),
		.single_rx_detect_hwtcl                   (0),
		.hip_hard_reset_hwtcl                     (1),
		.use_cvp_update_core_pof_hwtcl            (0),
		.pcie_inspector_hwtcl                     (0),
		.tlp_inspector_hwtcl                      (0),
		.tlp_inspector_use_signal_probe_hwtcl     (0),
		.tlp_insp_trg_dw0_hwtcl                   (2049),
		.tlp_insp_trg_dw1_hwtcl                   (0),
		.tlp_insp_trg_dw2_hwtcl                   (0),
		.tlp_insp_trg_dw3_hwtcl                   (0),
		.hwtcl_override_g2_txvod                  (1),
		.rpre_emph_a_val_hwtcl                    (9),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (16),
		.rpre_emph_d_val_hwtcl                    (13),
		.rpre_emph_e_val_hwtcl                    (5),
		.rvod_sel_a_val_hwtcl                     (42),
		.rvod_sel_b_val_hwtcl                     (38),
		.rvod_sel_c_val_hwtcl                     (38),
		.rvod_sel_d_val_hwtcl                     (43),
		.rvod_sel_e_val_hwtcl                     (15)
	) pcie (
		.coreclkout           (pcie_coreclkout_clk),                      //          coreclkout.clk
		.refclk               (pcie_refclk_clk),                          //              refclk.clk
		.npor                 (pcie_npor_npor),                           //                npor.npor
		.pin_perst            (pcie_npor_pin_perst),                      //                    .pin_perst
		.reset_status         (pcie_nreset_status_reset),                 //       nreset_status.reset_n
		.RxmAddress_0_o       (pcie_rxm_bar0_address),                    //            Rxm_BAR0.address
		.RxmRead_0_o          (pcie_rxm_bar0_read),                       //                    .read
		.RxmWaitRequest_0_i   (pcie_rxm_bar0_waitrequest),                //                    .waitrequest
		.RxmWrite_0_o         (pcie_rxm_bar0_write),                      //                    .write
		.RxmReadDataValid_0_i (pcie_rxm_bar0_readdatavalid),              //                    .readdatavalid
		.RxmReadData_0_i      (pcie_rxm_bar0_readdata),                   //                    .readdata
		.RxmWriteData_0_o     (pcie_rxm_bar0_writedata),                  //                    .writedata
		.RxmBurstCount_0_o    (pcie_rxm_bar0_burstcount),                 //                    .burstcount
		.RxmByteEnable_0_o    (pcie_rxm_bar0_byteenable),                 //                    .byteenable
		.RxmIrq_i             (pcie_rxmirq_irq),                          //              RxmIrq.irq
		.reconfig_to_xcvr     (reconfig_to_xcvr_reconfig_to_xcvr),        //    reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr   (reconfig_from_xcvr_reconfig_from_xcvr),    //  reconfig_from_xcvr.reconfig_from_xcvr
		.fixedclk_locked      (),                                         // reconfig_clk_locked.fixedclk_locked
		.rx_in0               (pcie_hip_serial_rx_in0),                   //          hip_serial.rx_in0
		.rx_in1               (pcie_hip_serial_rx_in1),                   //                    .rx_in1
		.rx_in2               (pcie_hip_serial_rx_in2),                   //                    .rx_in2
		.rx_in3               (pcie_hip_serial_rx_in3),                   //                    .rx_in3
		.rx_in4               (pcie_hip_serial_rx_in4),                   //                    .rx_in4
		.rx_in5               (pcie_hip_serial_rx_in5),                   //                    .rx_in5
		.rx_in6               (pcie_hip_serial_rx_in6),                   //                    .rx_in6
		.rx_in7               (pcie_hip_serial_rx_in7),                   //                    .rx_in7
		.tx_out0              (pcie_hip_serial_tx_out0),                  //                    .tx_out0
		.tx_out1              (pcie_hip_serial_tx_out1),                  //                    .tx_out1
		.tx_out2              (pcie_hip_serial_tx_out2),                  //                    .tx_out2
		.tx_out3              (pcie_hip_serial_tx_out3),                  //                    .tx_out3
		.tx_out4              (pcie_hip_serial_tx_out4),                  //                    .tx_out4
		.tx_out5              (pcie_hip_serial_tx_out5),                  //                    .tx_out5
		.tx_out6              (pcie_hip_serial_tx_out6),                  //                    .tx_out6
		.tx_out7              (pcie_hip_serial_tx_out7),                  //                    .tx_out7
		.sim_pipe_pclk_in     (),                                         //            hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate        (),                                         //                    .sim_pipe_rate
		.sim_ltssmstate       (),                                         //                    .sim_ltssmstate
		.eidleinfersel0       (),                                         //                    .eidleinfersel0
		.eidleinfersel1       (),                                         //                    .eidleinfersel1
		.eidleinfersel2       (),                                         //                    .eidleinfersel2
		.eidleinfersel3       (),                                         //                    .eidleinfersel3
		.eidleinfersel4       (),                                         //                    .eidleinfersel4
		.eidleinfersel5       (),                                         //                    .eidleinfersel5
		.eidleinfersel6       (),                                         //                    .eidleinfersel6
		.eidleinfersel7       (),                                         //                    .eidleinfersel7
		.powerdown0           (),                                         //                    .powerdown0
		.powerdown1           (),                                         //                    .powerdown1
		.powerdown2           (),                                         //                    .powerdown2
		.powerdown3           (),                                         //                    .powerdown3
		.powerdown4           (),                                         //                    .powerdown4
		.powerdown5           (),                                         //                    .powerdown5
		.powerdown6           (),                                         //                    .powerdown6
		.powerdown7           (),                                         //                    .powerdown7
		.rxpolarity0          (),                                         //                    .rxpolarity0
		.rxpolarity1          (),                                         //                    .rxpolarity1
		.rxpolarity2          (),                                         //                    .rxpolarity2
		.rxpolarity3          (),                                         //                    .rxpolarity3
		.rxpolarity4          (),                                         //                    .rxpolarity4
		.rxpolarity5          (),                                         //                    .rxpolarity5
		.rxpolarity6          (),                                         //                    .rxpolarity6
		.rxpolarity7          (),                                         //                    .rxpolarity7
		.txcompl0             (),                                         //                    .txcompl0
		.txcompl1             (),                                         //                    .txcompl1
		.txcompl2             (),                                         //                    .txcompl2
		.txcompl3             (),                                         //                    .txcompl3
		.txcompl4             (),                                         //                    .txcompl4
		.txcompl5             (),                                         //                    .txcompl5
		.txcompl6             (),                                         //                    .txcompl6
		.txcompl7             (),                                         //                    .txcompl7
		.txdata0              (),                                         //                    .txdata0
		.txdata1              (),                                         //                    .txdata1
		.txdata2              (),                                         //                    .txdata2
		.txdata3              (),                                         //                    .txdata3
		.txdata4              (),                                         //                    .txdata4
		.txdata5              (),                                         //                    .txdata5
		.txdata6              (),                                         //                    .txdata6
		.txdata7              (),                                         //                    .txdata7
		.txdatak0             (),                                         //                    .txdatak0
		.txdatak1             (),                                         //                    .txdatak1
		.txdatak2             (),                                         //                    .txdatak2
		.txdatak3             (),                                         //                    .txdatak3
		.txdatak4             (),                                         //                    .txdatak4
		.txdatak5             (),                                         //                    .txdatak5
		.txdatak6             (),                                         //                    .txdatak6
		.txdatak7             (),                                         //                    .txdatak7
		.txdetectrx0          (),                                         //                    .txdetectrx0
		.txdetectrx1          (),                                         //                    .txdetectrx1
		.txdetectrx2          (),                                         //                    .txdetectrx2
		.txdetectrx3          (),                                         //                    .txdetectrx3
		.txdetectrx4          (),                                         //                    .txdetectrx4
		.txdetectrx5          (),                                         //                    .txdetectrx5
		.txdetectrx6          (),                                         //                    .txdetectrx6
		.txdetectrx7          (),                                         //                    .txdetectrx7
		.txelecidle0          (),                                         //                    .txelecidle0
		.txelecidle1          (),                                         //                    .txelecidle1
		.txelecidle2          (),                                         //                    .txelecidle2
		.txelecidle3          (),                                         //                    .txelecidle3
		.txelecidle4          (),                                         //                    .txelecidle4
		.txelecidle5          (),                                         //                    .txelecidle5
		.txelecidle6          (),                                         //                    .txelecidle6
		.txelecidle7          (),                                         //                    .txelecidle7
		.txdeemph0            (),                                         //                    .txdeemph0
		.txdeemph1            (),                                         //                    .txdeemph1
		.txdeemph2            (),                                         //                    .txdeemph2
		.txdeemph3            (),                                         //                    .txdeemph3
		.txdeemph4            (),                                         //                    .txdeemph4
		.txdeemph5            (),                                         //                    .txdeemph5
		.txdeemph6            (),                                         //                    .txdeemph6
		.txdeemph7            (),                                         //                    .txdeemph7
		.txmargin0            (),                                         //                    .txmargin0
		.txmargin1            (),                                         //                    .txmargin1
		.txmargin2            (),                                         //                    .txmargin2
		.txmargin3            (),                                         //                    .txmargin3
		.txmargin4            (),                                         //                    .txmargin4
		.txmargin5            (),                                         //                    .txmargin5
		.txmargin6            (),                                         //                    .txmargin6
		.txmargin7            (),                                         //                    .txmargin7
		.txswing0             (),                                         //                    .txswing0
		.txswing1             (),                                         //                    .txswing1
		.txswing2             (),                                         //                    .txswing2
		.txswing3             (),                                         //                    .txswing3
		.txswing4             (),                                         //                    .txswing4
		.txswing5             (),                                         //                    .txswing5
		.txswing6             (),                                         //                    .txswing6
		.txswing7             (),                                         //                    .txswing7
		.phystatus0           (),                                         //                    .phystatus0
		.phystatus1           (),                                         //                    .phystatus1
		.phystatus2           (),                                         //                    .phystatus2
		.phystatus3           (),                                         //                    .phystatus3
		.phystatus4           (),                                         //                    .phystatus4
		.phystatus5           (),                                         //                    .phystatus5
		.phystatus6           (),                                         //                    .phystatus6
		.phystatus7           (),                                         //                    .phystatus7
		.rxdata0              (),                                         //                    .rxdata0
		.rxdata1              (),                                         //                    .rxdata1
		.rxdata2              (),                                         //                    .rxdata2
		.rxdata3              (),                                         //                    .rxdata3
		.rxdata4              (),                                         //                    .rxdata4
		.rxdata5              (),                                         //                    .rxdata5
		.rxdata6              (),                                         //                    .rxdata6
		.rxdata7              (),                                         //                    .rxdata7
		.rxdatak0             (),                                         //                    .rxdatak0
		.rxdatak1             (),                                         //                    .rxdatak1
		.rxdatak2             (),                                         //                    .rxdatak2
		.rxdatak3             (),                                         //                    .rxdatak3
		.rxdatak4             (),                                         //                    .rxdatak4
		.rxdatak5             (),                                         //                    .rxdatak5
		.rxdatak6             (),                                         //                    .rxdatak6
		.rxdatak7             (),                                         //                    .rxdatak7
		.rxelecidle0          (),                                         //                    .rxelecidle0
		.rxelecidle1          (),                                         //                    .rxelecidle1
		.rxelecidle2          (),                                         //                    .rxelecidle2
		.rxelecidle3          (),                                         //                    .rxelecidle3
		.rxelecidle4          (),                                         //                    .rxelecidle4
		.rxelecidle5          (),                                         //                    .rxelecidle5
		.rxelecidle6          (),                                         //                    .rxelecidle6
		.rxelecidle7          (),                                         //                    .rxelecidle7
		.rxstatus0            (),                                         //                    .rxstatus0
		.rxstatus1            (),                                         //                    .rxstatus1
		.rxstatus2            (),                                         //                    .rxstatus2
		.rxstatus3            (),                                         //                    .rxstatus3
		.rxstatus4            (),                                         //                    .rxstatus4
		.rxstatus5            (),                                         //                    .rxstatus5
		.rxstatus6            (),                                         //                    .rxstatus6
		.rxstatus7            (),                                         //                    .rxstatus7
		.rxvalid0             (),                                         //                    .rxvalid0
		.rxvalid1             (),                                         //                    .rxvalid1
		.rxvalid2             (),                                         //                    .rxvalid2
		.rxvalid3             (),                                         //                    .rxvalid3
		.rxvalid4             (),                                         //                    .rxvalid4
		.rxvalid5             (),                                         //                    .rxvalid5
		.rxvalid6             (),                                         //                    .rxvalid6
		.rxvalid7             (),                                         //                    .rxvalid7
		.test_in              (pcie_hip_ctrl_test_in),                    //            hip_ctrl.test_in
		.simu_mode_pipe       (pcie_hip_ctrl_simu_mode_pipe),             //                    .simu_mode_pipe
		.TxsChipSelect_i      (mm_interconnect_9_pcie_txs_chipselect),    //                 Txs.chipselect
		.TxsByteEnable_i      (mm_interconnect_9_pcie_txs_byteenable),    //                    .byteenable
		.TxsReadData_o        (mm_interconnect_9_pcie_txs_readdata),      //                    .readdata
		.TxsWriteData_i       (mm_interconnect_9_pcie_txs_writedata),     //                    .writedata
		.TxsRead_i            (mm_interconnect_9_pcie_txs_read),          //                    .read
		.TxsWrite_i           (mm_interconnect_9_pcie_txs_write),         //                    .write
		.TxsBurstCount_i      (mm_interconnect_9_pcie_txs_burstcount),    //                    .burstcount
		.TxsReadDataValid_o   (mm_interconnect_9_pcie_txs_readdatavalid), //                    .readdatavalid
		.TxsWaitRequest_o     (mm_interconnect_9_pcie_txs_waitrequest),   //                    .waitrequest
		.TxsAddress_i         (mm_interconnect_9_pcie_txs_address),       //                    .address
		.CraChipSelect_i      (mm_interconnect_2_pcie_cra_chipselect),    //                 Cra.chipselect
		.CraAddress_i         (mm_interconnect_2_pcie_cra_address),       //                    .address
		.CraByteEnable_i      (mm_interconnect_2_pcie_cra_byteenable),    //                    .byteenable
		.CraRead              (mm_interconnect_2_pcie_cra_read),          //                    .read
		.CraReadData_o        (mm_interconnect_2_pcie_cra_readdata),      //                    .readdata
		.CraWrite             (mm_interconnect_2_pcie_cra_write),         //                    .write
		.CraWriteData_i       (mm_interconnect_2_pcie_cra_writedata),     //                    .writedata
		.CraWaitRequest_o     (mm_interconnect_2_pcie_cra_waitrequest),   //                    .waitrequest
		.CraIrq_o             (),                                         //              CraIrq.irq
		.rxdataskip0          (1'b0),                                     //         (terminated)
		.rxdataskip1          (1'b0),                                     //         (terminated)
		.rxdataskip2          (1'b0),                                     //         (terminated)
		.rxdataskip3          (1'b0),                                     //         (terminated)
		.rxdataskip4          (1'b0),                                     //         (terminated)
		.rxdataskip5          (1'b0),                                     //         (terminated)
		.rxdataskip6          (1'b0),                                     //         (terminated)
		.rxdataskip7          (1'b0),                                     //         (terminated)
		.rxblkst0             (1'b0),                                     //         (terminated)
		.rxblkst1             (1'b0),                                     //         (terminated)
		.rxblkst2             (1'b0),                                     //         (terminated)
		.rxblkst3             (1'b0),                                     //         (terminated)
		.rxblkst4             (1'b0),                                     //         (terminated)
		.rxblkst5             (1'b0),                                     //         (terminated)
		.rxblkst6             (1'b0),                                     //         (terminated)
		.rxblkst7             (1'b0),                                     //         (terminated)
		.rxsynchd0            (2'b00),                                    //         (terminated)
		.rxsynchd1            (2'b00),                                    //         (terminated)
		.rxsynchd2            (2'b00),                                    //         (terminated)
		.rxsynchd3            (2'b00),                                    //         (terminated)
		.rxsynchd4            (2'b00),                                    //         (terminated)
		.rxsynchd5            (2'b00),                                    //         (terminated)
		.rxsynchd6            (2'b00),                                    //         (terminated)
		.rxsynchd7            (2'b00),                                    //         (terminated)
		.rxfreqlocked0        (1'b0),                                     //         (terminated)
		.rxfreqlocked1        (1'b0),                                     //         (terminated)
		.rxfreqlocked2        (1'b0),                                     //         (terminated)
		.rxfreqlocked3        (1'b0),                                     //         (terminated)
		.rxfreqlocked4        (1'b0),                                     //         (terminated)
		.rxfreqlocked5        (1'b0),                                     //         (terminated)
		.rxfreqlocked6        (1'b0),                                     //         (terminated)
		.rxfreqlocked7        (1'b0),                                     //         (terminated)
		.currentcoeff0        (),                                         //         (terminated)
		.currentcoeff1        (),                                         //         (terminated)
		.currentcoeff2        (),                                         //         (terminated)
		.currentcoeff3        (),                                         //         (terminated)
		.currentcoeff4        (),                                         //         (terminated)
		.currentcoeff5        (),                                         //         (terminated)
		.currentcoeff6        (),                                         //         (terminated)
		.currentcoeff7        (),                                         //         (terminated)
		.currentrxpreset0     (),                                         //         (terminated)
		.currentrxpreset1     (),                                         //         (terminated)
		.currentrxpreset2     (),                                         //         (terminated)
		.currentrxpreset3     (),                                         //         (terminated)
		.currentrxpreset4     (),                                         //         (terminated)
		.currentrxpreset5     (),                                         //         (terminated)
		.currentrxpreset6     (),                                         //         (terminated)
		.currentrxpreset7     (),                                         //         (terminated)
		.txsynchd0            (),                                         //         (terminated)
		.txsynchd1            (),                                         //         (terminated)
		.txsynchd2            (),                                         //         (terminated)
		.txsynchd3            (),                                         //         (terminated)
		.txsynchd4            (),                                         //         (terminated)
		.txsynchd5            (),                                         //         (terminated)
		.txsynchd6            (),                                         //         (terminated)
		.txsynchd7            (),                                         //         (terminated)
		.txblkst0             (),                                         //         (terminated)
		.txblkst1             (),                                         //         (terminated)
		.txblkst2             (),                                         //         (terminated)
		.txblkst3             (),                                         //         (terminated)
		.txblkst4             (),                                         //         (terminated)
		.txblkst5             (),                                         //         (terminated)
		.txblkst6             (),                                         //         (terminated)
		.txblkst7             ()                                          //         (terminated)
	);

	system_acl_iface_ddr3a ddr3a (
		.pll_ref_clk               (ddr3a_pll_ref_clk),                              //      pll_ref_clk.clk
		.global_reset_n            (~reset_controller_global_reset_out_reset),       //     global_reset.reset_n
		.soft_reset_n              (~reset_controller_global_reset_out_reset),       //       soft_reset.reset_n
		.afi_clk                   (ddr3a_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (),                                               //     afi_half_clk.clk
		.afi_reset_n               (),                                               //        afi_reset.reset_n
		.afi_reset_export_n        (),                                               // afi_reset_export.reset_n
		.mem_a                     (ddr3a_mem_a),                                    //           memory.mem_a
		.mem_ba                    (ddr3a_mem_ba),                                   //                 .mem_ba
		.mem_ck                    (ddr3a_mem_ck),                                   //                 .mem_ck
		.mem_ck_n                  (ddr3a_mem_ck_n),                                 //                 .mem_ck_n
		.mem_cke                   (ddr3a_mem_cke),                                  //                 .mem_cke
		.mem_cs_n                  (ddr3a_mem_cs_n),                                 //                 .mem_cs_n
		.mem_dm                    (ddr3a_mem_dm),                                   //                 .mem_dm
		.mem_ras_n                 (ddr3a_mem_ras_n),                                //                 .mem_ras_n
		.mem_cas_n                 (ddr3a_mem_cas_n),                                //                 .mem_cas_n
		.mem_we_n                  (ddr3a_mem_we_n),                                 //                 .mem_we_n
		.mem_reset_n               (ddr3a_mem_reset_n),                              //                 .mem_reset_n
		.mem_dq                    (ddr3a_mem_dq),                                   //                 .mem_dq
		.mem_dqs                   (ddr3a_mem_dqs),                                  //                 .mem_dqs
		.mem_dqs_n                 (ddr3a_mem_dqs_n),                                //                 .mem_dqs_n
		.mem_odt                   (ddr3a_mem_odt),                                  //                 .mem_odt
		.avl_ready                 (mm_interconnect_0_ddr3a_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_0_ddr3a_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_0_ddr3a_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_0_ddr3a_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_0_ddr3a_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_0_ddr3a_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_0_ddr3a_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_0_ddr3a_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_0_ddr3a_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_0_ddr3a_avl_burstcount),         //                 .burstcount
		.local_init_done           (ddr3a_status_local_init_done),                   //           status.local_init_done
		.local_cal_success         (ddr3a_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail            (ddr3a_status_local_cal_fail),                    //                 .local_cal_fail
		.oct_rzqin                 (octa_rzqin),                                     //              oct.rzqin
		.pll_mem_clk               (),                                               //      pll_sharing.pll_mem_clk
		.pll_write_clk             (),                                               //                 .pll_write_clk
		.pll_locked                (),                                               //                 .pll_locked
		.pll_write_clk_pre_phy_clk (),                                               //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (),                                               //                 .pll_addr_cmd_clk
		.pll_avl_clk               (),                                               //                 .pll_avl_clk
		.pll_config_clk            (),                                               //                 .pll_config_clk
		.pll_hr_clk                (),                                               //                 .pll_hr_clk
		.pll_p2c_read_clk          (),                                               //                 .pll_p2c_read_clk
		.pll_c2p_write_clk         ()                                                //                 .pll_c2p_write_clk
	);

	system_acl_iface_ddr3b ddr3b (
		.pll_ref_clk               (ddr3b_pll_ref_clk),                              //      pll_ref_clk.clk
		.global_reset_n            (~reset_controller_global_reset_out_reset),       //     global_reset.reset_n
		.soft_reset_n              (~reset_controller_global_reset_out_reset),       //       soft_reset.reset_n
		.afi_clk                   (ddr3b_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (),                                               //     afi_half_clk.clk
		.afi_reset_n               (),                                               //        afi_reset.reset_n
		.afi_reset_export_n        (),                                               // afi_reset_export.reset_n
		.mem_a                     (ddr3b_mem_a),                                    //           memory.mem_a
		.mem_ba                    (ddr3b_mem_ba),                                   //                 .mem_ba
		.mem_ck                    (ddr3b_mem_ck),                                   //                 .mem_ck
		.mem_ck_n                  (ddr3b_mem_ck_n),                                 //                 .mem_ck_n
		.mem_cke                   (ddr3b_mem_cke),                                  //                 .mem_cke
		.mem_cs_n                  (ddr3b_mem_cs_n),                                 //                 .mem_cs_n
		.mem_dm                    (ddr3b_mem_dm),                                   //                 .mem_dm
		.mem_ras_n                 (ddr3b_mem_ras_n),                                //                 .mem_ras_n
		.mem_cas_n                 (ddr3b_mem_cas_n),                                //                 .mem_cas_n
		.mem_we_n                  (ddr3b_mem_we_n),                                 //                 .mem_we_n
		.mem_reset_n               (ddr3b_mem_reset_n),                              //                 .mem_reset_n
		.mem_dq                    (ddr3b_mem_dq),                                   //                 .mem_dq
		.mem_dqs                   (ddr3b_mem_dqs),                                  //                 .mem_dqs
		.mem_dqs_n                 (ddr3b_mem_dqs_n),                                //                 .mem_dqs_n
		.mem_odt                   (ddr3b_mem_odt),                                  //                 .mem_odt
		.avl_ready                 (mm_interconnect_1_ddr3b_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_1_ddr3b_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_1_ddr3b_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_1_ddr3b_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_1_ddr3b_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_1_ddr3b_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_1_ddr3b_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_1_ddr3b_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_1_ddr3b_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_1_ddr3b_avl_burstcount),         //                 .burstcount
		.local_init_done           (ddr3b_status_local_init_done),                   //           status.local_init_done
		.local_cal_success         (ddr3b_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail            (ddr3b_status_local_cal_fail),                    //                 .local_cal_fail
		.oct_rzqin                 (octb_rzqin),                                     //              oct.rzqin
		.pll_mem_clk               (),                                               //      pll_sharing.pll_mem_clk
		.pll_write_clk             (),                                               //                 .pll_write_clk
		.pll_locked                (),                                               //                 .pll_locked
		.pll_write_clk_pre_phy_clk (),                                               //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (),                                               //                 .pll_addr_cmd_clk
		.pll_avl_clk               (),                                               //                 .pll_avl_clk
		.pll_config_clk            (),                                               //                 .pll_config_clk
		.pll_hr_clk                (),                                               //                 .pll_hr_clk
		.pll_p2c_read_clk          (),                                               //                 .pll_p2c_read_clk
		.pll_c2p_write_clk         ()                                                //                 .pll_c2p_write_clk
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (512),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (31),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pipe_stage_ddr3a_dimm (
		.clk              (ddr3a_afi_clk_clk),                       //   clk.clk
		.reset            (reset_controller_ddr3a_reset_out_reset),  // reset.reset
		.s0_waitrequest   (pipe_stage_ddr3a_iface_m0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (pipe_stage_ddr3a_iface_m0_readdata),      //      .readdata
		.s0_readdatavalid (pipe_stage_ddr3a_iface_m0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (pipe_stage_ddr3a_iface_m0_burstcount),    //      .burstcount
		.s0_writedata     (pipe_stage_ddr3a_iface_m0_writedata),     //      .writedata
		.s0_address       (pipe_stage_ddr3a_iface_m0_address),       //      .address
		.s0_write         (pipe_stage_ddr3a_iface_m0_write),         //      .write
		.s0_read          (pipe_stage_ddr3a_iface_m0_read),          //      .read
		.s0_byteenable    (pipe_stage_ddr3a_iface_m0_byteenable),    //      .byteenable
		.s0_debugaccess   (pipe_stage_ddr3a_iface_m0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pipe_stage_ddr3a_dimm_m0_waitrequest),    //    m0.waitrequest
		.m0_readdata      (pipe_stage_ddr3a_dimm_m0_readdata),       //      .readdata
		.m0_readdatavalid (pipe_stage_ddr3a_dimm_m0_readdatavalid),  //      .readdatavalid
		.m0_burstcount    (pipe_stage_ddr3a_dimm_m0_burstcount),     //      .burstcount
		.m0_writedata     (pipe_stage_ddr3a_dimm_m0_writedata),      //      .writedata
		.m0_address       (pipe_stage_ddr3a_dimm_m0_address),        //      .address
		.m0_write         (pipe_stage_ddr3a_dimm_m0_write),          //      .write
		.m0_read          (pipe_stage_ddr3a_dimm_m0_read),           //      .read
		.m0_byteenable    (pipe_stage_ddr3a_dimm_m0_byteenable),     //      .byteenable
		.m0_debugaccess   (pipe_stage_ddr3a_dimm_m0_debugaccess),    //      .debugaccess
		.s0_response      (),                                        // (terminated)
		.m0_response      (2'b00)                                    // (terminated)
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (512),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (20),
		.BURSTCOUNT_WIDTH    (5),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) clock_cross_dma_to_pcie (
		.m0_clk           (pcie_coreclkout_clk),                                        //   m0_clk.clk
		.m0_reset         (reset_controller_pcie_reset_out_reset),                      // m0_reset.reset
		.s0_clk           (ddr3a_afi_clk_clk),                                          //   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset),                             // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_3_clock_cross_dma_to_pcie_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_3_clock_cross_dma_to_pcie_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_3_clock_cross_dma_to_pcie_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_3_clock_cross_dma_to_pcie_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_3_clock_cross_dma_to_pcie_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_3_clock_cross_dma_to_pcie_s0_address),       //         .address
		.s0_write         (mm_interconnect_3_clock_cross_dma_to_pcie_s0_write),         //         .write
		.s0_read          (mm_interconnect_3_clock_cross_dma_to_pcie_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_3_clock_cross_dma_to_pcie_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_3_clock_cross_dma_to_pcie_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_cross_dma_to_pcie_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_cross_dma_to_pcie_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_cross_dma_to_pcie_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_cross_dma_to_pcie_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_cross_dma_to_pcie_m0_writedata),                       //         .writedata
		.m0_address       (clock_cross_dma_to_pcie_m0_address),                         //         .address
		.m0_write         (clock_cross_dma_to_pcie_m0_write),                           //         .write
		.m0_read          (clock_cross_dma_to_pcie_m0_read),                            //         .read
		.m0_byteenable    (clock_cross_dma_to_pcie_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_cross_dma_to_pcie_m0_debugaccess)                      //         .debugaccess
	);

	system_acl_iface_temperature_pll temperature_pll (
		.refclk   (config_clk_clk),                          //  refclk.clk
		.rst      (reset_controller_global_reset_out_reset), //   reset.reset
		.outclk_0 (temperature_pll_outclk0_clk),             // outclk0.clk
		.locked   ()                                         //  locked.export
	);

	temperature temperature_0 (
		.clk                 (temperature_pll_outclk0_clk),                     //       clk.clk
		.resetn              (~rst_controller_001_reset_out_reset),             // clk_reset.reset_n
		.slave_address       (mm_interconnect_2_temperature_0_s_address),       //         s.address
		.slave_writedata     (mm_interconnect_2_temperature_0_s_writedata),     //          .writedata
		.slave_read          (mm_interconnect_2_temperature_0_s_read),          //          .read
		.slave_write         (mm_interconnect_2_temperature_0_s_write),         //          .write
		.slave_byteenable    (mm_interconnect_2_temperature_0_s_byteenable),    //          .byteenable
		.slave_waitrequest   (mm_interconnect_2_temperature_0_s_waitrequest),   //          .waitrequest
		.slave_readdata      (mm_interconnect_2_temperature_0_s_readdata),      //          .readdata
		.slave_readdatavalid (mm_interconnect_2_temperature_0_s_readdatavalid)  //          .readdatavalid
	);

	system_acl_iface_acl_kernel_clk acl_kernel_clk (
		.pll_refclk_clk           (kernel_pll_refclk_clk),                               //        pll_refclk.clk
		.clk_clk                  (config_clk_clk),                                      //               clk.clk
		.reset_reset_n            (~reset_controller_global_reset_out_reset),            //             reset.reset_n
		.ctrl_waitrequest         (mm_interconnect_2_acl_kernel_clk_ctrl_waitrequest),   //              ctrl.waitrequest
		.ctrl_readdata            (mm_interconnect_2_acl_kernel_clk_ctrl_readdata),      //                  .readdata
		.ctrl_readdatavalid       (mm_interconnect_2_acl_kernel_clk_ctrl_readdatavalid), //                  .readdatavalid
		.ctrl_burstcount          (mm_interconnect_2_acl_kernel_clk_ctrl_burstcount),    //                  .burstcount
		.ctrl_writedata           (mm_interconnect_2_acl_kernel_clk_ctrl_writedata),     //                  .writedata
		.ctrl_address             (mm_interconnect_2_acl_kernel_clk_ctrl_address),       //                  .address
		.ctrl_write               (mm_interconnect_2_acl_kernel_clk_ctrl_write),         //                  .write
		.ctrl_read                (mm_interconnect_2_acl_kernel_clk_ctrl_read),          //                  .read
		.ctrl_byteenable          (mm_interconnect_2_acl_kernel_clk_ctrl_byteenable),    //                  .byteenable
		.ctrl_debugaccess         (mm_interconnect_2_acl_kernel_clk_ctrl_debugaccess),   //                  .debugaccess
		.kernel_clk_clk           (kernel_clk_clk),                                      //        kernel_clk.clk
		.kernel_clk2x_clk         (kernel_clk2x_clk),                                    //      kernel_clk2x.clk
		.kernel_pll_locked_export ()                                                     // kernel_pll_locked.export
	);

	system_acl_iface_kernel_interface kernel_interface (
		.clk_clk                    (pcie_coreclkout_clk),                                           //                    clk.clk
		.reset_reset_n              (~reset_controller_pcie_reset_out_reset),                        //                  reset.reset_n
		.kernel_cntrl_waitrequest   (mm_interconnect_2_kernel_interface_kernel_cntrl_waitrequest),   //           kernel_cntrl.waitrequest
		.kernel_cntrl_readdata      (mm_interconnect_2_kernel_interface_kernel_cntrl_readdata),      //                       .readdata
		.kernel_cntrl_readdatavalid (mm_interconnect_2_kernel_interface_kernel_cntrl_readdatavalid), //                       .readdatavalid
		.kernel_cntrl_burstcount    (mm_interconnect_2_kernel_interface_kernel_cntrl_burstcount),    //                       .burstcount
		.kernel_cntrl_writedata     (mm_interconnect_2_kernel_interface_kernel_cntrl_writedata),     //                       .writedata
		.kernel_cntrl_address       (mm_interconnect_2_kernel_interface_kernel_cntrl_address),       //                       .address
		.kernel_cntrl_write         (mm_interconnect_2_kernel_interface_kernel_cntrl_write),         //                       .write
		.kernel_cntrl_read          (mm_interconnect_2_kernel_interface_kernel_cntrl_read),          //                       .read
		.kernel_cntrl_byteenable    (mm_interconnect_2_kernel_interface_kernel_cntrl_byteenable),    //                       .byteenable
		.kernel_cntrl_debugaccess   (mm_interconnect_2_kernel_interface_kernel_cntrl_debugaccess),   //                       .debugaccess
		.kernel_clk_clk             (kernel_clk_clk),                                                //             kernel_clk.clk
		.kernel_cra_waitrequest     (kernel_cra_waitrequest),                                        //             kernel_cra.waitrequest
		.kernel_cra_readdata        (kernel_cra_readdata),                                           //                       .readdata
		.kernel_cra_readdatavalid   (kernel_cra_readdatavalid),                                      //                       .readdatavalid
		.kernel_cra_burstcount      (kernel_cra_burstcount),                                         //                       .burstcount
		.kernel_cra_writedata       (kernel_cra_writedata),                                          //                       .writedata
		.kernel_cra_address         (kernel_cra_address),                                            //                       .address
		.kernel_cra_write           (kernel_cra_write),                                              //                       .write
		.kernel_cra_read            (kernel_cra_read),                                               //                       .read
		.kernel_cra_byteenable      (kernel_cra_byteenable),                                         //                       .byteenable
		.kernel_cra_debugaccess     (kernel_cra_debugaccess),                                        //                       .debugaccess
		.sw_reset_in_reset          (reset_controller_pcie_reset_out_reset),                         //            sw_reset_in.reset
		.kernel_reset_reset_n       (kernel_reset_reset_n),                                          //           kernel_reset.reset_n
		.sw_reset_export_reset_n    (kernel_interface_sw_reset_export_reset),                        //        sw_reset_export.reset_n
		.acl_bsp_memorg_kernel_mode (acl_internal_memorg_kernel_mode),                               //  acl_bsp_memorg_kernel.mode
		.acl_bsp_memorg_host_mode   (kernel_interface_acl_bsp_memorg_host_mode),                     //    acl_bsp_memorg_host.mode
		.kernel_irq_from_kernel_irq (kernel_irq_irq),                                                // kernel_irq_from_kernel.irq
		.kernel_irq_to_host_irq     (irq_synchronizer_receiver_irq)                                  //     kernel_irq_to_host.irq
	);

	system_acl_iface_dma_0 dma_0 (
		.dma_irq_irq            (irq_synchronizer_001_receiver_irq),              //  dma_irq.irq
		.reset_reset_n          (~rst_controller_002_reset_out_reset),            //    reset.reset_n
		.clk_clk                (ddr3a_afi_clk_clk),                              //      clk.clk
		.m_waitrequest          (dma_0_m_waitrequest),                            //        m.waitrequest
		.m_readdata             (dma_0_m_readdata),                               //         .readdata
		.m_readdatavalid        (dma_0_m_readdatavalid),                          //         .readdatavalid
		.m_burstcount           (dma_0_m_burstcount),                             //         .burstcount
		.m_writedata            (dma_0_m_writedata),                              //         .writedata
		.m_address              (dma_0_m_address),                                //         .address
		.m_write                (dma_0_m_write),                                  //         .write
		.m_read                 (dma_0_m_read),                                   //         .read
		.m_byteenable           (dma_0_m_byteenable),                             //         .byteenable
		.m_debugaccess          (dma_0_m_debugaccess),                            //         .debugaccess
		.csr_waitrequest        (mm_interconnect_2_dma_0_csr_waitrequest),        //      csr.waitrequest
		.csr_readdata           (mm_interconnect_2_dma_0_csr_readdata),           //         .readdata
		.csr_readdatavalid      (mm_interconnect_2_dma_0_csr_readdatavalid),      //         .readdatavalid
		.csr_burstcount         (mm_interconnect_2_dma_0_csr_burstcount),         //         .burstcount
		.csr_writedata          (mm_interconnect_2_dma_0_csr_writedata),          //         .writedata
		.csr_address            (mm_interconnect_2_dma_0_csr_address),            //         .address
		.csr_write              (mm_interconnect_2_dma_0_csr_write),              //         .write
		.csr_read               (mm_interconnect_2_dma_0_csr_read),               //         .read
		.csr_byteenable         (mm_interconnect_2_dma_0_csr_byteenable),         //         .byteenable
		.csr_debugaccess        (mm_interconnect_2_dma_0_csr_debugaccess),        //         .debugaccess
		.s_nondma_address       (mm_interconnect_2_dma_0_s_nondma_address),       // s_nondma.address
		.s_nondma_read          (mm_interconnect_2_dma_0_s_nondma_read),          //         .read
		.s_nondma_readdata      (mm_interconnect_2_dma_0_s_nondma_readdata),      //         .readdata
		.s_nondma_write         (mm_interconnect_2_dma_0_s_nondma_write),         //         .write
		.s_nondma_writedata     (mm_interconnect_2_dma_0_s_nondma_writedata),     //         .writedata
		.s_nondma_readdatavalid (mm_interconnect_2_dma_0_s_nondma_readdatavalid), //         .readdatavalid
		.s_nondma_waitrequest   (mm_interconnect_2_dma_0_s_nondma_waitrequest),   //         .waitrequest
		.s_nondma_byteenable    (mm_interconnect_2_dma_0_s_nondma_byteenable),    //         .byteenable
		.s_nondma_burstcount    (mm_interconnect_2_dma_0_s_nondma_burstcount)     //         .burstcount
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (18),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pipe_stage_host_ctrl (
		.clk              (pcie_coreclkout_clk),                                     //   clk.clk
		.reset            (reset_controller_pcie_reset_out_reset),                   // reset.reset
		.s0_waitrequest   (mm_interconnect_8_pipe_stage_host_ctrl_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_8_pipe_stage_host_ctrl_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_8_pipe_stage_host_ctrl_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_8_pipe_stage_host_ctrl_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_8_pipe_stage_host_ctrl_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_8_pipe_stage_host_ctrl_s0_address),       //      .address
		.s0_write         (mm_interconnect_8_pipe_stage_host_ctrl_s0_write),         //      .write
		.s0_read          (mm_interconnect_8_pipe_stage_host_ctrl_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_8_pipe_stage_host_ctrl_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_8_pipe_stage_host_ctrl_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pipe_stage_host_ctrl_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (pipe_stage_host_ctrl_m0_readdata),                        //      .readdata
		.m0_readdatavalid (pipe_stage_host_ctrl_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (pipe_stage_host_ctrl_m0_burstcount),                      //      .burstcount
		.m0_writedata     (pipe_stage_host_ctrl_m0_writedata),                       //      .writedata
		.m0_address       (pipe_stage_host_ctrl_m0_address),                         //      .address
		.m0_write         (pipe_stage_host_ctrl_m0_write),                           //      .write
		.m0_read          (pipe_stage_host_ctrl_m0_read),                            //      .read
		.m0_byteenable    (pipe_stage_host_ctrl_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (pipe_stage_host_ctrl_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                        // (terminated)
		.m0_response      (2'b00)                                                    // (terminated)
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (512),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (31),
		.BURSTCOUNT_WIDTH    (5),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (512),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) clock_cross_kernel_mem_0 (
		.m0_clk           (ddr3a_afi_clk_clk),                         //   m0_clk.clk
		.m0_reset         (rst_controller_003_reset_out_reset),        // m0_reset.reset
		.s0_clk           (kernel_clk_clk),                            //   s0_clk.clk
		.s0_reset         (~kernel_reset_reset_n),                     // s0_reset.reset
		.s0_waitrequest   (kernel_mem0_waitrequest),                   //       s0.waitrequest
		.s0_readdata      (kernel_mem0_readdata),                      //         .readdata
		.s0_readdatavalid (kernel_mem0_readdatavalid),                 //         .readdatavalid
		.s0_burstcount    (kernel_mem0_burstcount),                    //         .burstcount
		.s0_writedata     (kernel_mem0_writedata),                     //         .writedata
		.s0_address       (kernel_mem0_address),                       //         .address
		.s0_write         (kernel_mem0_write),                         //         .write
		.s0_read          (kernel_mem0_read),                          //         .read
		.s0_byteenable    (kernel_mem0_byteenable),                    //         .byteenable
		.s0_debugaccess   (kernel_mem0_debugaccess),                   //         .debugaccess
		.m0_waitrequest   (clock_cross_kernel_mem_0_m0_waitrequest),   //       m0.waitrequest
		.m0_readdata      (clock_cross_kernel_mem_0_m0_readdata),      //         .readdata
		.m0_readdatavalid (clock_cross_kernel_mem_0_m0_readdatavalid), //         .readdatavalid
		.m0_burstcount    (clock_cross_kernel_mem_0_m0_burstcount),    //         .burstcount
		.m0_writedata     (clock_cross_kernel_mem_0_m0_writedata),     //         .writedata
		.m0_address       (clock_cross_kernel_mem_0_m0_address),       //         .address
		.m0_write         (clock_cross_kernel_mem_0_m0_write),         //         .write
		.m0_read          (clock_cross_kernel_mem_0_m0_read),          //         .read
		.m0_byteenable    (clock_cross_kernel_mem_0_m0_byteenable),    //         .byteenable
		.m0_debugaccess   (clock_cross_kernel_mem_0_m0_debugaccess)    //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (512),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (31),
		.BURSTCOUNT_WIDTH    (5),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (512),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) clock_cross_kernel_mem_1 (
		.m0_clk           (ddr3b_afi_clk_clk),                         //   m0_clk.clk
		.m0_reset         (rst_controller_004_reset_out_reset),        // m0_reset.reset
		.s0_clk           (kernel_clk_clk),                            //   s0_clk.clk
		.s0_reset         (~kernel_reset_reset_n),                     // s0_reset.reset
		.s0_waitrequest   (kernel_mem1_waitrequest),                   //       s0.waitrequest
		.s0_readdata      (kernel_mem1_readdata),                      //         .readdata
		.s0_readdatavalid (kernel_mem1_readdatavalid),                 //         .readdatavalid
		.s0_burstcount    (kernel_mem1_burstcount),                    //         .burstcount
		.s0_writedata     (kernel_mem1_writedata),                     //         .writedata
		.s0_address       (kernel_mem1_address),                       //         .address
		.s0_write         (kernel_mem1_write),                         //         .write
		.s0_read          (kernel_mem1_read),                          //         .read
		.s0_byteenable    (kernel_mem1_byteenable),                    //         .byteenable
		.s0_debugaccess   (kernel_mem1_debugaccess),                   //         .debugaccess
		.m0_waitrequest   (clock_cross_kernel_mem_1_m0_waitrequest),   //       m0.waitrequest
		.m0_readdata      (clock_cross_kernel_mem_1_m0_readdata),      //         .readdata
		.m0_readdatavalid (clock_cross_kernel_mem_1_m0_readdatavalid), //         .readdatavalid
		.m0_burstcount    (clock_cross_kernel_mem_1_m0_burstcount),    //         .burstcount
		.m0_writedata     (clock_cross_kernel_mem_1_m0_writedata),     //         .writedata
		.m0_address       (clock_cross_kernel_mem_1_m0_address),       //         .address
		.m0_write         (clock_cross_kernel_mem_1_m0_write),         //         .write
		.m0_read          (clock_cross_kernel_mem_1_m0_read),          //         .read
		.m0_byteenable    (clock_cross_kernel_mem_1_m0_byteenable),    //         .byteenable
		.m0_debugaccess   (clock_cross_kernel_mem_1_m0_debugaccess)    //         .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (512),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (31),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pipe_stage_ddr3a_iface (
		.clk              (ddr3a_afi_clk_clk),                                         //   clk.clk
		.reset            (reset_controller_ddr3a_reset_out_reset),                    // reset.reset
		.s0_waitrequest   (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_address),       //      .address
		.s0_write         (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_write),         //      .write
		.s0_read          (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pipe_stage_ddr3a_iface_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (pipe_stage_ddr3a_iface_m0_readdata),                        //      .readdata
		.m0_readdatavalid (pipe_stage_ddr3a_iface_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (pipe_stage_ddr3a_iface_m0_burstcount),                      //      .burstcount
		.m0_writedata     (pipe_stage_ddr3a_iface_m0_writedata),                       //      .writedata
		.m0_address       (pipe_stage_ddr3a_iface_m0_address),                         //      .address
		.m0_write         (pipe_stage_ddr3a_iface_m0_write),                           //      .write
		.m0_read          (pipe_stage_ddr3a_iface_m0_read),                            //      .read
		.m0_byteenable    (pipe_stage_ddr3a_iface_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (pipe_stage_ddr3a_iface_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                          // (terminated)
		.m0_response      (2'b00)                                                      // (terminated)
	);

	system_acl_iface_em_pc_0 #(
		.EMPC_AV_BURSTCOUNT_WIDTH (1),
		.EMPC_AV_DATA_WIDTH       (512),
		.EMPC_AV_POW2_DATA_WIDTH  (512),
		.EMPC_AV_ADDRESS_WIDTH    (25),
		.EMPC_AV_SYMBOL_WIDTH     (8),
		.EMPC_COUNT_WIDTH         (32)
	) em_pc_0 (
		.avl_in_address             (mm_interconnect_5_em_pc_0_avl_in_address),            //      avl_in.address
		.avl_in_byteenable          (mm_interconnect_5_em_pc_0_avl_in_byteenable),         //            .byteenable
		.avl_in_burstcount          (mm_interconnect_5_em_pc_0_avl_in_burstcount),         //            .burstcount
		.avl_in_beginbursttransfer  (mm_interconnect_5_em_pc_0_avl_in_beginbursttransfer), //            .beginbursttransfer
		.avl_in_waitrequest         (mm_interconnect_5_em_pc_0_avl_in_waitrequest),        //            .waitrequest
		.avl_in_write               (mm_interconnect_5_em_pc_0_avl_in_write),              //            .write
		.avl_in_read                (mm_interconnect_5_em_pc_0_avl_in_read),               //            .read
		.avl_in_readdatavalid       (mm_interconnect_5_em_pc_0_avl_in_readdatavalid),      //            .readdatavalid
		.avl_in_writedata           (mm_interconnect_5_em_pc_0_avl_in_writedata),          //            .writedata
		.avl_in_readdata            (mm_interconnect_5_em_pc_0_avl_in_readdata),           //            .readdata
		.avl_out_address            (em_pc_0_avl_out_address),                             //     avl_out.address
		.avl_out_byteenable         (em_pc_0_avl_out_byteenable),                          //            .byteenable
		.avl_out_burstcount         (em_pc_0_avl_out_burstcount),                          //            .burstcount
		.avl_out_beginbursttransfer (em_pc_0_avl_out_beginbursttransfer),                  //            .beginbursttransfer
		.avl_out_waitrequest        (em_pc_0_avl_out_waitrequest),                         //            .waitrequest
		.avl_out_write              (em_pc_0_avl_out_write),                               //            .write
		.avl_out_read               (em_pc_0_avl_out_read),                                //            .read
		.avl_out_readdatavalid      (em_pc_0_avl_out_readdatavalid),                       //            .readdatavalid
		.avl_out_writedata          (em_pc_0_avl_out_writedata),                           //            .writedata
		.avl_out_readdata           (em_pc_0_avl_out_readdata),                            //            .readdata
		.avl_clk                    (ddr3a_afi_clk_clk),                                   //     avl_clk.clk
		.avl_reset_n                (~reset_controller_ddr3a_reset_out_reset),             // avl_reset_n.reset_n
		.em_csr_waitrequest         (mm_interconnect_2_em_pc_0_em_csr_waitrequest),        //      em_csr.waitrequest
		.em_csr_readdata            (mm_interconnect_2_em_pc_0_em_csr_readdata),           //            .readdata
		.em_csr_readdatavalid       (mm_interconnect_2_em_pc_0_em_csr_readdatavalid),      //            .readdatavalid
		.em_csr_burstcount          (mm_interconnect_2_em_pc_0_em_csr_burstcount),         //            .burstcount
		.em_csr_writedata           (mm_interconnect_2_em_pc_0_em_csr_writedata),          //            .writedata
		.em_csr_address             (mm_interconnect_2_em_pc_0_em_csr_address),            //            .address
		.em_csr_write               (mm_interconnect_2_em_pc_0_em_csr_write),              //            .write
		.em_csr_read                (mm_interconnect_2_em_pc_0_em_csr_read),               //            .read
		.em_csr_byteenable          (mm_interconnect_2_em_pc_0_em_csr_byteenable),         //            .byteenable
		.em_csr_debugaccess         (mm_interconnect_2_em_pc_0_em_csr_debugaccess)         //            .debugaccess
	);

	system_acl_iface_em_pc_0 #(
		.EMPC_AV_BURSTCOUNT_WIDTH (1),
		.EMPC_AV_DATA_WIDTH       (512),
		.EMPC_AV_POW2_DATA_WIDTH  (512),
		.EMPC_AV_ADDRESS_WIDTH    (25),
		.EMPC_AV_SYMBOL_WIDTH     (8),
		.EMPC_COUNT_WIDTH         (32)
	) em_pc_1 (
		.avl_in_address             (mm_interconnect_7_em_pc_1_avl_in_address),            //      avl_in.address
		.avl_in_byteenable          (mm_interconnect_7_em_pc_1_avl_in_byteenable),         //            .byteenable
		.avl_in_burstcount          (mm_interconnect_7_em_pc_1_avl_in_burstcount),         //            .burstcount
		.avl_in_beginbursttransfer  (mm_interconnect_7_em_pc_1_avl_in_beginbursttransfer), //            .beginbursttransfer
		.avl_in_waitrequest         (mm_interconnect_7_em_pc_1_avl_in_waitrequest),        //            .waitrequest
		.avl_in_write               (mm_interconnect_7_em_pc_1_avl_in_write),              //            .write
		.avl_in_read                (mm_interconnect_7_em_pc_1_avl_in_read),               //            .read
		.avl_in_readdatavalid       (mm_interconnect_7_em_pc_1_avl_in_readdatavalid),      //            .readdatavalid
		.avl_in_writedata           (mm_interconnect_7_em_pc_1_avl_in_writedata),          //            .writedata
		.avl_in_readdata            (mm_interconnect_7_em_pc_1_avl_in_readdata),           //            .readdata
		.avl_out_address            (em_pc_1_avl_out_address),                             //     avl_out.address
		.avl_out_byteenable         (em_pc_1_avl_out_byteenable),                          //            .byteenable
		.avl_out_burstcount         (em_pc_1_avl_out_burstcount),                          //            .burstcount
		.avl_out_beginbursttransfer (em_pc_1_avl_out_beginbursttransfer),                  //            .beginbursttransfer
		.avl_out_waitrequest        (em_pc_1_avl_out_waitrequest),                         //            .waitrequest
		.avl_out_write              (em_pc_1_avl_out_write),                               //            .write
		.avl_out_read               (em_pc_1_avl_out_read),                                //            .read
		.avl_out_readdatavalid      (em_pc_1_avl_out_readdatavalid),                       //            .readdatavalid
		.avl_out_writedata          (em_pc_1_avl_out_writedata),                           //            .writedata
		.avl_out_readdata           (em_pc_1_avl_out_readdata),                            //            .readdata
		.avl_clk                    (ddr3b_afi_clk_clk),                                   //     avl_clk.clk
		.avl_reset_n                (~reset_controller_ddr3b_reset_out_reset),             // avl_reset_n.reset_n
		.em_csr_waitrequest         (mm_interconnect_2_em_pc_1_em_csr_waitrequest),        //      em_csr.waitrequest
		.em_csr_readdata            (mm_interconnect_2_em_pc_1_em_csr_readdata),           //            .readdata
		.em_csr_readdatavalid       (mm_interconnect_2_em_pc_1_em_csr_readdatavalid),      //            .readdatavalid
		.em_csr_burstcount          (mm_interconnect_2_em_pc_1_em_csr_burstcount),         //            .burstcount
		.em_csr_writedata           (mm_interconnect_2_em_pc_1_em_csr_writedata),          //            .writedata
		.em_csr_address             (mm_interconnect_2_em_pc_1_em_csr_address),            //            .address
		.em_csr_write               (mm_interconnect_2_em_pc_1_em_csr_write),              //            .write
		.em_csr_read                (mm_interconnect_2_em_pc_1_em_csr_read),               //            .read
		.em_csr_byteenable          (mm_interconnect_2_em_pc_1_em_csr_byteenable),         //            .byteenable
		.em_csr_debugaccess         (mm_interconnect_2_em_pc_1_em_csr_debugaccess)         //            .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (512),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (31),
		.BURSTCOUNT_WIDTH    (5),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) clock_cross_dma_to_ddr3b (
		.m0_clk           (ddr3b_afi_clk_clk),                                            //   m0_clk.clk
		.m0_reset         (reset_controller_ddr3b_reset_out_reset),                       // m0_reset.reset
		.s0_clk           (ddr3a_afi_clk_clk),                                            //   s0_clk.clk
		.s0_reset         (reset_controller_ddr3a_reset_out_reset),                       // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_address),       //         .address
		.s0_write         (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_write),         //         .write
		.s0_read          (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_cross_dma_to_ddr3b_m0_waitrequest),                      //       m0.waitrequest
		.m0_readdata      (clock_cross_dma_to_ddr3b_m0_readdata),                         //         .readdata
		.m0_readdatavalid (clock_cross_dma_to_ddr3b_m0_readdatavalid),                    //         .readdatavalid
		.m0_burstcount    (clock_cross_dma_to_ddr3b_m0_burstcount),                       //         .burstcount
		.m0_writedata     (clock_cross_dma_to_ddr3b_m0_writedata),                        //         .writedata
		.m0_address       (clock_cross_dma_to_ddr3b_m0_address),                          //         .address
		.m0_write         (clock_cross_dma_to_ddr3b_m0_write),                            //         .write
		.m0_read          (clock_cross_dma_to_ddr3b_m0_read),                             //         .read
		.m0_byteenable    (clock_cross_dma_to_ddr3b_m0_byteenable),                       //         .byteenable
		.m0_debugaccess   (clock_cross_dma_to_ddr3b_m0_debugaccess)                       //         .debugaccess
	);

	system_acl_iface_acl_memory_bank_divider_0 acl_memory_bank_divider_0 (
		.clk_clk                  (ddr3a_afi_clk_clk),                                                //                 clk.clk
		.reset_reset_n            (~rst_controller_002_reset_out_reset),                              //               reset.reset_n
		.kernel_clk_clk           (kernel_clk_clk),                                                   //          kernel_clk.clk
		.kernel_reset_reset_n     (kernel_reset_reset_n),                                             //        kernel_reset.reset_n
		.acl_bsp_snoop_data       (acl_internal_snoop_data),                                          //       acl_bsp_snoop.data
		.acl_bsp_snoop_valid      (acl_internal_snoop_valid),                                         //                    .valid
		.acl_bsp_snoop_ready      (acl_internal_snoop_ready),                                         //                    .ready
		.s_read                   (mm_interconnect_3_acl_memory_bank_divider_0_s_read),               //                   s.read
		.s_readdata               (mm_interconnect_3_acl_memory_bank_divider_0_s_readdata),           //                    .readdata
		.s_readdatavalid          (mm_interconnect_3_acl_memory_bank_divider_0_s_readdatavalid),      //                    .readdatavalid
		.s_write                  (mm_interconnect_3_acl_memory_bank_divider_0_s_write),              //                    .write
		.s_writedata              (mm_interconnect_3_acl_memory_bank_divider_0_s_writedata),          //                    .writedata
		.s_burstcount             (mm_interconnect_3_acl_memory_bank_divider_0_s_burstcount),         //                    .burstcount
		.s_beginbursttransfer     (mm_interconnect_3_acl_memory_bank_divider_0_s_beginbursttransfer), //                    .beginbursttransfer
		.s_byteenable             (mm_interconnect_3_acl_memory_bank_divider_0_s_byteenable),         //                    .byteenable
		.s_address                (mm_interconnect_3_acl_memory_bank_divider_0_s_address),            //                    .address
		.s_waitrequest            (mm_interconnect_3_acl_memory_bank_divider_0_s_waitrequest),        //                    .waitrequest
		.acl_bsp_memorg_host_mode (kernel_interface_acl_bsp_memorg_host_mode),                        // acl_bsp_memorg_host.mode
		.bank1_address            (acl_memory_bank_divider_0_bank1_address),                          //               bank1.address
		.bank1_writedata          (acl_memory_bank_divider_0_bank1_writedata),                        //                    .writedata
		.bank1_read               (acl_memory_bank_divider_0_bank1_read),                             //                    .read
		.bank1_write              (acl_memory_bank_divider_0_bank1_write),                            //                    .write
		.bank1_burstcount         (acl_memory_bank_divider_0_bank1_burstcount),                       //                    .burstcount
		.bank1_byteenable         (acl_memory_bank_divider_0_bank1_byteenable),                       //                    .byteenable
		.bank1_waitrequest        (acl_memory_bank_divider_0_bank1_waitrequest),                      //                    .waitrequest
		.bank1_readdata           (acl_memory_bank_divider_0_bank1_readdata),                         //                    .readdata
		.bank1_readdatavalid      (acl_memory_bank_divider_0_bank1_readdatavalid),                    //                    .readdatavalid
		.bank2_address            (acl_memory_bank_divider_0_bank2_address),                          //               bank2.address
		.bank2_writedata          (acl_memory_bank_divider_0_bank2_writedata),                        //                    .writedata
		.bank2_read               (acl_memory_bank_divider_0_bank2_read),                             //                    .read
		.bank2_write              (acl_memory_bank_divider_0_bank2_write),                            //                    .write
		.bank2_burstcount         (acl_memory_bank_divider_0_bank2_burstcount),                       //                    .burstcount
		.bank2_byteenable         (acl_memory_bank_divider_0_bank2_byteenable),                       //                    .byteenable
		.bank2_waitrequest        (acl_memory_bank_divider_0_bank2_waitrequest),                      //                    .waitrequest
		.bank2_readdata           (acl_memory_bank_divider_0_bank2_readdata),                         //                    .readdata
		.bank2_readdatavalid      (acl_memory_bank_divider_0_bank2_readdatavalid)                     //                    .readdatavalid
	);

	sw_reset #(
		.WIDTH             (8),
		.LOG2_RESET_CYCLES (10)
	) por_reset_counter (
		.clk               (config_clk_clk),                      //       clk.clk
		.resetn            (~rst_controller_005_reset_out_reset), // clk_reset.reset_n
		.slave_write       (),                                    //         s.write
		.slave_writedata   (),                                    //          .writedata
		.slave_byteenable  (),                                    //          .byteenable
		.slave_read        (),                                    //          .read
		.slave_readdata    (),                                    //          .readdata
		.slave_waitrequest (),                                    //          .waitrequest
		.sw_reset_n_out    (pcie_npor_out_reset_n)                //  sw_reset.reset_n
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_controller_pcie (
		.reset_in0      (reset_controller_global_reset_out_reset), // reset_in0.reset
		.clk            (pcie_coreclkout_clk),                     //       clk.clk
		.reset_out      (reset_controller_pcie_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                        // (terminated)
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_in1      (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_controller_ddr3b (
		.reset_in0      (reset_controller_global_reset_out_reset), // reset_in0.reset
		.clk            (ddr3b_afi_clk_clk),                       //       clk.clk
		.reset_out      (reset_controller_ddr3b_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                        // (terminated)
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_in1      (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_controller_ddr3a (
		.reset_in0      (reset_controller_global_reset_out_reset), // reset_in0.reset
		.clk            (ddr3a_afi_clk_clk),                       //       clk.clk
		.reset_out      (reset_controller_ddr3a_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                        // (terminated)
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_in1      (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_controller_global (
		.reset_in0      (~pcie_npor_out_reset_n),                  // reset_in0.reset
		.reset_in1      (~pcie_nreset_status_reset),               // reset_in1.reset
		.clk            (config_clk_clk),                          //       clk.clk
		.reset_out      (reset_controller_global_reset_out_reset), // reset_out.reset
		.reset_req      (),                                        // (terminated)
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	uniphy_status #(
		.WIDTH       (32),
		.NUM_UNIPHYS (2)
	) uniphy_status_0 (
		.clk                      (pcie_coreclkout_clk),                          //           clk.clk
		.resetn                   (~rst_controller_006_reset_out_reset),          //     clk_reset.reset_n
		.mem0_local_init_done     (ddr3a_status_local_init_done),                 //   mem0_status.local_init_done
		.mem0_local_cal_success   (ddr3a_status_local_cal_success),               //              .local_cal_success
		.mem0_local_cal_fail      (ddr3a_status_local_cal_fail),                  //              .local_cal_fail
		.mem1_local_init_done     (ddr3b_status_local_init_done),                 //   mem1_status.local_init_done
		.mem1_local_cal_success   (ddr3b_status_local_cal_success),               //              .local_cal_success
		.mem1_local_cal_fail      (ddr3b_status_local_cal_fail),                  //              .local_cal_fail
		.export_local_init_done   (),                                             // status_export.local_init_done
		.export_local_cal_success (),                                             //              .local_cal_success
		.export_local_cal_fail    (),                                             //              .local_cal_fail
		.slave_read               (mm_interconnect_2_uniphy_status_0_s_read),     //             s.read
		.slave_readdata           (mm_interconnect_2_uniphy_status_0_s_readdata)  //              .readdata
	);

	version_id #(
		.WIDTH      (32),
		.VERSION_ID (-1597521440)
	) version_id_0 (
		.clk            (pcie_coreclkout_clk),                       //       clk.clk
		.resetn         (~rst_controller_006_reset_out_reset),       // clk_reset.reset_n
		.slave_read     (mm_interconnect_2_version_id_0_s_read),     //         s.read
		.slave_readdata (mm_interconnect_2_version_id_0_s_readdata)  //          .readdata
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (512),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (31),
		.BURSTCOUNT_WIDTH  (5),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pipe_stage_ddr3b_iface (
		.clk              (ddr3b_afi_clk_clk),                                          //   clk.clk
		.reset            (reset_controller_ddr3b_reset_out_reset),                     // reset.reset
		.s0_waitrequest   (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_address),       //      .address
		.s0_write         (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_write),         //      .write
		.s0_read          (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pipe_stage_ddr3b_iface_m0_waitrequest),                      //    m0.waitrequest
		.m0_readdata      (pipe_stage_ddr3b_iface_m0_readdata),                         //      .readdata
		.m0_readdatavalid (pipe_stage_ddr3b_iface_m0_readdatavalid),                    //      .readdatavalid
		.m0_burstcount    (pipe_stage_ddr3b_iface_m0_burstcount),                       //      .burstcount
		.m0_writedata     (pipe_stage_ddr3b_iface_m0_writedata),                        //      .writedata
		.m0_address       (pipe_stage_ddr3b_iface_m0_address),                          //      .address
		.m0_write         (pipe_stage_ddr3b_iface_m0_write),                            //      .write
		.m0_read          (pipe_stage_ddr3b_iface_m0_read),                             //      .read
		.m0_byteenable    (pipe_stage_ddr3b_iface_m0_byteenable),                       //      .byteenable
		.m0_debugaccess   (pipe_stage_ddr3b_iface_m0_debugaccess),                      //      .debugaccess
		.s0_response      (),                                                           // (terminated)
		.m0_response      (2'b00)                                                       // (terminated)
	);

	system_acl_iface_mm_interconnect_0 mm_interconnect_0 (
		.ddr3a_afi_clk_clk                                       (ddr3a_afi_clk_clk),                              //                                     ddr3a_afi_clk.clk
		.ddr3a_avl_translator_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                 //  ddr3a_avl_translator_reset_reset_bridge_in_reset.reset
		.ddr3a_soft_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                 //            ddr3a_soft_reset_reset_bridge_in_reset.reset
		.pipe_stage_ddr3a_dimm_reset_reset_bridge_in_reset_reset (reset_controller_ddr3a_reset_out_reset),         // pipe_stage_ddr3a_dimm_reset_reset_bridge_in_reset.reset
		.pipe_stage_ddr3a_dimm_m0_address                        (pipe_stage_ddr3a_dimm_m0_address),               //                          pipe_stage_ddr3a_dimm_m0.address
		.pipe_stage_ddr3a_dimm_m0_waitrequest                    (pipe_stage_ddr3a_dimm_m0_waitrequest),           //                                                  .waitrequest
		.pipe_stage_ddr3a_dimm_m0_burstcount                     (pipe_stage_ddr3a_dimm_m0_burstcount),            //                                                  .burstcount
		.pipe_stage_ddr3a_dimm_m0_byteenable                     (pipe_stage_ddr3a_dimm_m0_byteenable),            //                                                  .byteenable
		.pipe_stage_ddr3a_dimm_m0_read                           (pipe_stage_ddr3a_dimm_m0_read),                  //                                                  .read
		.pipe_stage_ddr3a_dimm_m0_readdata                       (pipe_stage_ddr3a_dimm_m0_readdata),              //                                                  .readdata
		.pipe_stage_ddr3a_dimm_m0_readdatavalid                  (pipe_stage_ddr3a_dimm_m0_readdatavalid),         //                                                  .readdatavalid
		.pipe_stage_ddr3a_dimm_m0_write                          (pipe_stage_ddr3a_dimm_m0_write),                 //                                                  .write
		.pipe_stage_ddr3a_dimm_m0_writedata                      (pipe_stage_ddr3a_dimm_m0_writedata),             //                                                  .writedata
		.pipe_stage_ddr3a_dimm_m0_debugaccess                    (pipe_stage_ddr3a_dimm_m0_debugaccess),           //                                                  .debugaccess
		.ddr3a_avl_address                                       (mm_interconnect_0_ddr3a_avl_address),            //                                         ddr3a_avl.address
		.ddr3a_avl_write                                         (mm_interconnect_0_ddr3a_avl_write),              //                                                  .write
		.ddr3a_avl_read                                          (mm_interconnect_0_ddr3a_avl_read),               //                                                  .read
		.ddr3a_avl_readdata                                      (mm_interconnect_0_ddr3a_avl_readdata),           //                                                  .readdata
		.ddr3a_avl_writedata                                     (mm_interconnect_0_ddr3a_avl_writedata),          //                                                  .writedata
		.ddr3a_avl_beginbursttransfer                            (mm_interconnect_0_ddr3a_avl_beginbursttransfer), //                                                  .beginbursttransfer
		.ddr3a_avl_burstcount                                    (mm_interconnect_0_ddr3a_avl_burstcount),         //                                                  .burstcount
		.ddr3a_avl_byteenable                                    (mm_interconnect_0_ddr3a_avl_byteenable),         //                                                  .byteenable
		.ddr3a_avl_readdatavalid                                 (mm_interconnect_0_ddr3a_avl_readdatavalid),      //                                                  .readdatavalid
		.ddr3a_avl_waitrequest                                   (~mm_interconnect_0_ddr3a_avl_waitrequest)        //                                                  .waitrequest
	);

	system_acl_iface_mm_interconnect_1 mm_interconnect_1 (
		.ddr3b_afi_clk_clk                                       (ddr3b_afi_clk_clk),                              //                                     ddr3b_afi_clk.clk
		.ddr3b_avl_translator_reset_reset_bridge_in_reset_reset  (rst_controller_007_reset_out_reset),             //  ddr3b_avl_translator_reset_reset_bridge_in_reset.reset
		.ddr3b_soft_reset_reset_bridge_in_reset_reset            (rst_controller_007_reset_out_reset),             //            ddr3b_soft_reset_reset_bridge_in_reset.reset
		.pipe_stage_ddr3b_dimm_reset_reset_bridge_in_reset_reset (reset_controller_ddr3b_reset_out_reset),         // pipe_stage_ddr3b_dimm_reset_reset_bridge_in_reset.reset
		.pipe_stage_ddr3b_dimm_m0_address                        (pipe_stage_ddr3b_dimm_m0_address),               //                          pipe_stage_ddr3b_dimm_m0.address
		.pipe_stage_ddr3b_dimm_m0_waitrequest                    (pipe_stage_ddr3b_dimm_m0_waitrequest),           //                                                  .waitrequest
		.pipe_stage_ddr3b_dimm_m0_burstcount                     (pipe_stage_ddr3b_dimm_m0_burstcount),            //                                                  .burstcount
		.pipe_stage_ddr3b_dimm_m0_byteenable                     (pipe_stage_ddr3b_dimm_m0_byteenable),            //                                                  .byteenable
		.pipe_stage_ddr3b_dimm_m0_read                           (pipe_stage_ddr3b_dimm_m0_read),                  //                                                  .read
		.pipe_stage_ddr3b_dimm_m0_readdata                       (pipe_stage_ddr3b_dimm_m0_readdata),              //                                                  .readdata
		.pipe_stage_ddr3b_dimm_m0_readdatavalid                  (pipe_stage_ddr3b_dimm_m0_readdatavalid),         //                                                  .readdatavalid
		.pipe_stage_ddr3b_dimm_m0_write                          (pipe_stage_ddr3b_dimm_m0_write),                 //                                                  .write
		.pipe_stage_ddr3b_dimm_m0_writedata                      (pipe_stage_ddr3b_dimm_m0_writedata),             //                                                  .writedata
		.pipe_stage_ddr3b_dimm_m0_debugaccess                    (pipe_stage_ddr3b_dimm_m0_debugaccess),           //                                                  .debugaccess
		.ddr3b_avl_address                                       (mm_interconnect_1_ddr3b_avl_address),            //                                         ddr3b_avl.address
		.ddr3b_avl_write                                         (mm_interconnect_1_ddr3b_avl_write),              //                                                  .write
		.ddr3b_avl_read                                          (mm_interconnect_1_ddr3b_avl_read),               //                                                  .read
		.ddr3b_avl_readdata                                      (mm_interconnect_1_ddr3b_avl_readdata),           //                                                  .readdata
		.ddr3b_avl_writedata                                     (mm_interconnect_1_ddr3b_avl_writedata),          //                                                  .writedata
		.ddr3b_avl_beginbursttransfer                            (mm_interconnect_1_ddr3b_avl_beginbursttransfer), //                                                  .beginbursttransfer
		.ddr3b_avl_burstcount                                    (mm_interconnect_1_ddr3b_avl_burstcount),         //                                                  .burstcount
		.ddr3b_avl_byteenable                                    (mm_interconnect_1_ddr3b_avl_byteenable),         //                                                  .byteenable
		.ddr3b_avl_readdatavalid                                 (mm_interconnect_1_ddr3b_avl_readdatavalid),      //                                                  .readdatavalid
		.ddr3b_avl_waitrequest                                   (~mm_interconnect_1_ddr3b_avl_waitrequest)        //                                                  .waitrequest
	);

	system_acl_iface_mm_interconnect_2 mm_interconnect_2 (
		.config_clk_out_clk_clk                                      (config_clk_clk),                                                //                                    config_clk_out_clk.clk
		.ddr3a_afi_clk_clk                                           (ddr3a_afi_clk_clk),                                             //                                         ddr3a_afi_clk.clk
		.ddr3b_afi_clk_clk                                           (ddr3b_afi_clk_clk),                                             //                                         ddr3b_afi_clk.clk
		.pcie_coreclkout_clk                                         (pcie_coreclkout_clk),                                           //                                       pcie_coreclkout.clk
		.temperature_pll_outclk0_clk                                 (temperature_pll_outclk0_clk),                                   //                               temperature_pll_outclk0.clk
		.acl_kernel_clk_reset_reset_bridge_in_reset_reset            (reset_controller_global_reset_out_reset),                       //            acl_kernel_clk_reset_reset_bridge_in_reset.reset
		.dma_0_reset_reset_bridge_in_reset_reset                     (rst_controller_002_reset_out_reset),                            //                     dma_0_reset_reset_bridge_in_reset.reset
		.em_pc_0_avl_reset_n_reset_bridge_in_reset_reset             (reset_controller_ddr3a_reset_out_reset),                        //             em_pc_0_avl_reset_n_reset_bridge_in_reset.reset
		.em_pc_0_em_csr_translator_reset_reset_bridge_in_reset_reset (reset_controller_ddr3a_reset_out_reset),                        // em_pc_0_em_csr_translator_reset_reset_bridge_in_reset.reset
		.em_pc_1_avl_reset_n_reset_bridge_in_reset_reset             (reset_controller_ddr3b_reset_out_reset),                        //             em_pc_1_avl_reset_n_reset_bridge_in_reset.reset
		.em_pc_1_em_csr_translator_reset_reset_bridge_in_reset_reset (reset_controller_ddr3b_reset_out_reset),                        // em_pc_1_em_csr_translator_reset_reset_bridge_in_reset.reset
		.pcie_Cra_translator_reset_reset_bridge_in_reset_reset       (rst_controller_008_reset_out_reset),                            //       pcie_Cra_translator_reset_reset_bridge_in_reset.reset
		.pipe_stage_host_ctrl_reset_reset_bridge_in_reset_reset      (reset_controller_pcie_reset_out_reset),                         //      pipe_stage_host_ctrl_reset_reset_bridge_in_reset.reset
		.temperature_0_clk_reset_reset_bridge_in_reset_reset         (rst_controller_001_reset_out_reset),                            //         temperature_0_clk_reset_reset_bridge_in_reset.reset
		.uniphy_status_0_clk_reset_reset_bridge_in_reset_reset       (rst_controller_006_reset_out_reset),                            //       uniphy_status_0_clk_reset_reset_bridge_in_reset.reset
		.pipe_stage_host_ctrl_m0_address                             (pipe_stage_host_ctrl_m0_address),                               //                               pipe_stage_host_ctrl_m0.address
		.pipe_stage_host_ctrl_m0_waitrequest                         (pipe_stage_host_ctrl_m0_waitrequest),                           //                                                      .waitrequest
		.pipe_stage_host_ctrl_m0_burstcount                          (pipe_stage_host_ctrl_m0_burstcount),                            //                                                      .burstcount
		.pipe_stage_host_ctrl_m0_byteenable                          (pipe_stage_host_ctrl_m0_byteenable),                            //                                                      .byteenable
		.pipe_stage_host_ctrl_m0_read                                (pipe_stage_host_ctrl_m0_read),                                  //                                                      .read
		.pipe_stage_host_ctrl_m0_readdata                            (pipe_stage_host_ctrl_m0_readdata),                              //                                                      .readdata
		.pipe_stage_host_ctrl_m0_readdatavalid                       (pipe_stage_host_ctrl_m0_readdatavalid),                         //                                                      .readdatavalid
		.pipe_stage_host_ctrl_m0_write                               (pipe_stage_host_ctrl_m0_write),                                 //                                                      .write
		.pipe_stage_host_ctrl_m0_writedata                           (pipe_stage_host_ctrl_m0_writedata),                             //                                                      .writedata
		.pipe_stage_host_ctrl_m0_debugaccess                         (pipe_stage_host_ctrl_m0_debugaccess),                           //                                                      .debugaccess
		.acl_kernel_clk_ctrl_address                                 (mm_interconnect_2_acl_kernel_clk_ctrl_address),                 //                                   acl_kernel_clk_ctrl.address
		.acl_kernel_clk_ctrl_write                                   (mm_interconnect_2_acl_kernel_clk_ctrl_write),                   //                                                      .write
		.acl_kernel_clk_ctrl_read                                    (mm_interconnect_2_acl_kernel_clk_ctrl_read),                    //                                                      .read
		.acl_kernel_clk_ctrl_readdata                                (mm_interconnect_2_acl_kernel_clk_ctrl_readdata),                //                                                      .readdata
		.acl_kernel_clk_ctrl_writedata                               (mm_interconnect_2_acl_kernel_clk_ctrl_writedata),               //                                                      .writedata
		.acl_kernel_clk_ctrl_burstcount                              (mm_interconnect_2_acl_kernel_clk_ctrl_burstcount),              //                                                      .burstcount
		.acl_kernel_clk_ctrl_byteenable                              (mm_interconnect_2_acl_kernel_clk_ctrl_byteenable),              //                                                      .byteenable
		.acl_kernel_clk_ctrl_readdatavalid                           (mm_interconnect_2_acl_kernel_clk_ctrl_readdatavalid),           //                                                      .readdatavalid
		.acl_kernel_clk_ctrl_waitrequest                             (mm_interconnect_2_acl_kernel_clk_ctrl_waitrequest),             //                                                      .waitrequest
		.acl_kernel_clk_ctrl_debugaccess                             (mm_interconnect_2_acl_kernel_clk_ctrl_debugaccess),             //                                                      .debugaccess
		.dma_0_csr_address                                           (mm_interconnect_2_dma_0_csr_address),                           //                                             dma_0_csr.address
		.dma_0_csr_write                                             (mm_interconnect_2_dma_0_csr_write),                             //                                                      .write
		.dma_0_csr_read                                              (mm_interconnect_2_dma_0_csr_read),                              //                                                      .read
		.dma_0_csr_readdata                                          (mm_interconnect_2_dma_0_csr_readdata),                          //                                                      .readdata
		.dma_0_csr_writedata                                         (mm_interconnect_2_dma_0_csr_writedata),                         //                                                      .writedata
		.dma_0_csr_burstcount                                        (mm_interconnect_2_dma_0_csr_burstcount),                        //                                                      .burstcount
		.dma_0_csr_byteenable                                        (mm_interconnect_2_dma_0_csr_byteenable),                        //                                                      .byteenable
		.dma_0_csr_readdatavalid                                     (mm_interconnect_2_dma_0_csr_readdatavalid),                     //                                                      .readdatavalid
		.dma_0_csr_waitrequest                                       (mm_interconnect_2_dma_0_csr_waitrequest),                       //                                                      .waitrequest
		.dma_0_csr_debugaccess                                       (mm_interconnect_2_dma_0_csr_debugaccess),                       //                                                      .debugaccess
		.dma_0_s_nondma_address                                      (mm_interconnect_2_dma_0_s_nondma_address),                      //                                        dma_0_s_nondma.address
		.dma_0_s_nondma_write                                        (mm_interconnect_2_dma_0_s_nondma_write),                        //                                                      .write
		.dma_0_s_nondma_read                                         (mm_interconnect_2_dma_0_s_nondma_read),                         //                                                      .read
		.dma_0_s_nondma_readdata                                     (mm_interconnect_2_dma_0_s_nondma_readdata),                     //                                                      .readdata
		.dma_0_s_nondma_writedata                                    (mm_interconnect_2_dma_0_s_nondma_writedata),                    //                                                      .writedata
		.dma_0_s_nondma_burstcount                                   (mm_interconnect_2_dma_0_s_nondma_burstcount),                   //                                                      .burstcount
		.dma_0_s_nondma_byteenable                                   (mm_interconnect_2_dma_0_s_nondma_byteenable),                   //                                                      .byteenable
		.dma_0_s_nondma_readdatavalid                                (mm_interconnect_2_dma_0_s_nondma_readdatavalid),                //                                                      .readdatavalid
		.dma_0_s_nondma_waitrequest                                  (mm_interconnect_2_dma_0_s_nondma_waitrequest),                  //                                                      .waitrequest
		.em_pc_0_em_csr_address                                      (mm_interconnect_2_em_pc_0_em_csr_address),                      //                                        em_pc_0_em_csr.address
		.em_pc_0_em_csr_write                                        (mm_interconnect_2_em_pc_0_em_csr_write),                        //                                                      .write
		.em_pc_0_em_csr_read                                         (mm_interconnect_2_em_pc_0_em_csr_read),                         //                                                      .read
		.em_pc_0_em_csr_readdata                                     (mm_interconnect_2_em_pc_0_em_csr_readdata),                     //                                                      .readdata
		.em_pc_0_em_csr_writedata                                    (mm_interconnect_2_em_pc_0_em_csr_writedata),                    //                                                      .writedata
		.em_pc_0_em_csr_burstcount                                   (mm_interconnect_2_em_pc_0_em_csr_burstcount),                   //                                                      .burstcount
		.em_pc_0_em_csr_byteenable                                   (mm_interconnect_2_em_pc_0_em_csr_byteenable),                   //                                                      .byteenable
		.em_pc_0_em_csr_readdatavalid                                (mm_interconnect_2_em_pc_0_em_csr_readdatavalid),                //                                                      .readdatavalid
		.em_pc_0_em_csr_waitrequest                                  (mm_interconnect_2_em_pc_0_em_csr_waitrequest),                  //                                                      .waitrequest
		.em_pc_0_em_csr_debugaccess                                  (mm_interconnect_2_em_pc_0_em_csr_debugaccess),                  //                                                      .debugaccess
		.em_pc_1_em_csr_address                                      (mm_interconnect_2_em_pc_1_em_csr_address),                      //                                        em_pc_1_em_csr.address
		.em_pc_1_em_csr_write                                        (mm_interconnect_2_em_pc_1_em_csr_write),                        //                                                      .write
		.em_pc_1_em_csr_read                                         (mm_interconnect_2_em_pc_1_em_csr_read),                         //                                                      .read
		.em_pc_1_em_csr_readdata                                     (mm_interconnect_2_em_pc_1_em_csr_readdata),                     //                                                      .readdata
		.em_pc_1_em_csr_writedata                                    (mm_interconnect_2_em_pc_1_em_csr_writedata),                    //                                                      .writedata
		.em_pc_1_em_csr_burstcount                                   (mm_interconnect_2_em_pc_1_em_csr_burstcount),                   //                                                      .burstcount
		.em_pc_1_em_csr_byteenable                                   (mm_interconnect_2_em_pc_1_em_csr_byteenable),                   //                                                      .byteenable
		.em_pc_1_em_csr_readdatavalid                                (mm_interconnect_2_em_pc_1_em_csr_readdatavalid),                //                                                      .readdatavalid
		.em_pc_1_em_csr_waitrequest                                  (mm_interconnect_2_em_pc_1_em_csr_waitrequest),                  //                                                      .waitrequest
		.em_pc_1_em_csr_debugaccess                                  (mm_interconnect_2_em_pc_1_em_csr_debugaccess),                  //                                                      .debugaccess
		.kernel_interface_kernel_cntrl_address                       (mm_interconnect_2_kernel_interface_kernel_cntrl_address),       //                         kernel_interface_kernel_cntrl.address
		.kernel_interface_kernel_cntrl_write                         (mm_interconnect_2_kernel_interface_kernel_cntrl_write),         //                                                      .write
		.kernel_interface_kernel_cntrl_read                          (mm_interconnect_2_kernel_interface_kernel_cntrl_read),          //                                                      .read
		.kernel_interface_kernel_cntrl_readdata                      (mm_interconnect_2_kernel_interface_kernel_cntrl_readdata),      //                                                      .readdata
		.kernel_interface_kernel_cntrl_writedata                     (mm_interconnect_2_kernel_interface_kernel_cntrl_writedata),     //                                                      .writedata
		.kernel_interface_kernel_cntrl_burstcount                    (mm_interconnect_2_kernel_interface_kernel_cntrl_burstcount),    //                                                      .burstcount
		.kernel_interface_kernel_cntrl_byteenable                    (mm_interconnect_2_kernel_interface_kernel_cntrl_byteenable),    //                                                      .byteenable
		.kernel_interface_kernel_cntrl_readdatavalid                 (mm_interconnect_2_kernel_interface_kernel_cntrl_readdatavalid), //                                                      .readdatavalid
		.kernel_interface_kernel_cntrl_waitrequest                   (mm_interconnect_2_kernel_interface_kernel_cntrl_waitrequest),   //                                                      .waitrequest
		.kernel_interface_kernel_cntrl_debugaccess                   (mm_interconnect_2_kernel_interface_kernel_cntrl_debugaccess),   //                                                      .debugaccess
		.pcie_Cra_address                                            (mm_interconnect_2_pcie_cra_address),                            //                                              pcie_Cra.address
		.pcie_Cra_write                                              (mm_interconnect_2_pcie_cra_write),                              //                                                      .write
		.pcie_Cra_read                                               (mm_interconnect_2_pcie_cra_read),                               //                                                      .read
		.pcie_Cra_readdata                                           (mm_interconnect_2_pcie_cra_readdata),                           //                                                      .readdata
		.pcie_Cra_writedata                                          (mm_interconnect_2_pcie_cra_writedata),                          //                                                      .writedata
		.pcie_Cra_byteenable                                         (mm_interconnect_2_pcie_cra_byteenable),                         //                                                      .byteenable
		.pcie_Cra_waitrequest                                        (mm_interconnect_2_pcie_cra_waitrequest),                        //                                                      .waitrequest
		.pcie_Cra_chipselect                                         (mm_interconnect_2_pcie_cra_chipselect),                         //                                                      .chipselect
		.temperature_0_s_address                                     (mm_interconnect_2_temperature_0_s_address),                     //                                       temperature_0_s.address
		.temperature_0_s_write                                       (mm_interconnect_2_temperature_0_s_write),                       //                                                      .write
		.temperature_0_s_read                                        (mm_interconnect_2_temperature_0_s_read),                        //                                                      .read
		.temperature_0_s_readdata                                    (mm_interconnect_2_temperature_0_s_readdata),                    //                                                      .readdata
		.temperature_0_s_writedata                                   (mm_interconnect_2_temperature_0_s_writedata),                   //                                                      .writedata
		.temperature_0_s_byteenable                                  (mm_interconnect_2_temperature_0_s_byteenable),                  //                                                      .byteenable
		.temperature_0_s_readdatavalid                               (mm_interconnect_2_temperature_0_s_readdatavalid),               //                                                      .readdatavalid
		.temperature_0_s_waitrequest                                 (mm_interconnect_2_temperature_0_s_waitrequest),                 //                                                      .waitrequest
		.uniphy_status_0_s_read                                      (mm_interconnect_2_uniphy_status_0_s_read),                      //                                     uniphy_status_0_s.read
		.uniphy_status_0_s_readdata                                  (mm_interconnect_2_uniphy_status_0_s_readdata),                  //                                                      .readdata
		.version_id_0_s_read                                         (mm_interconnect_2_version_id_0_s_read),                         //                                        version_id_0_s.read
		.version_id_0_s_readdata                                     (mm_interconnect_2_version_id_0_s_readdata)                      //                                                      .readdata
	);

	system_acl_iface_mm_interconnect_3 mm_interconnect_3 (
		.ddr3a_afi_clk_clk                                            (ddr3a_afi_clk_clk),                                                //                                          ddr3a_afi_clk.clk
		.clock_cross_dma_to_pcie_s0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                   // clock_cross_dma_to_pcie_s0_reset_reset_bridge_in_reset.reset
		.dma_0_reset_reset_bridge_in_reset_reset                      (rst_controller_002_reset_out_reset),                               //                      dma_0_reset_reset_bridge_in_reset.reset
		.dma_0_m_address                                              (dma_0_m_address),                                                  //                                                dma_0_m.address
		.dma_0_m_waitrequest                                          (dma_0_m_waitrequest),                                              //                                                       .waitrequest
		.dma_0_m_burstcount                                           (dma_0_m_burstcount),                                               //                                                       .burstcount
		.dma_0_m_byteenable                                           (dma_0_m_byteenable),                                               //                                                       .byteenable
		.dma_0_m_read                                                 (dma_0_m_read),                                                     //                                                       .read
		.dma_0_m_readdata                                             (dma_0_m_readdata),                                                 //                                                       .readdata
		.dma_0_m_readdatavalid                                        (dma_0_m_readdatavalid),                                            //                                                       .readdatavalid
		.dma_0_m_write                                                (dma_0_m_write),                                                    //                                                       .write
		.dma_0_m_writedata                                            (dma_0_m_writedata),                                                //                                                       .writedata
		.dma_0_m_debugaccess                                          (dma_0_m_debugaccess),                                              //                                                       .debugaccess
		.acl_memory_bank_divider_0_s_address                          (mm_interconnect_3_acl_memory_bank_divider_0_s_address),            //                            acl_memory_bank_divider_0_s.address
		.acl_memory_bank_divider_0_s_write                            (mm_interconnect_3_acl_memory_bank_divider_0_s_write),              //                                                       .write
		.acl_memory_bank_divider_0_s_read                             (mm_interconnect_3_acl_memory_bank_divider_0_s_read),               //                                                       .read
		.acl_memory_bank_divider_0_s_readdata                         (mm_interconnect_3_acl_memory_bank_divider_0_s_readdata),           //                                                       .readdata
		.acl_memory_bank_divider_0_s_writedata                        (mm_interconnect_3_acl_memory_bank_divider_0_s_writedata),          //                                                       .writedata
		.acl_memory_bank_divider_0_s_beginbursttransfer               (mm_interconnect_3_acl_memory_bank_divider_0_s_beginbursttransfer), //                                                       .beginbursttransfer
		.acl_memory_bank_divider_0_s_burstcount                       (mm_interconnect_3_acl_memory_bank_divider_0_s_burstcount),         //                                                       .burstcount
		.acl_memory_bank_divider_0_s_byteenable                       (mm_interconnect_3_acl_memory_bank_divider_0_s_byteenable),         //                                                       .byteenable
		.acl_memory_bank_divider_0_s_readdatavalid                    (mm_interconnect_3_acl_memory_bank_divider_0_s_readdatavalid),      //                                                       .readdatavalid
		.acl_memory_bank_divider_0_s_waitrequest                      (mm_interconnect_3_acl_memory_bank_divider_0_s_waitrequest),        //                                                       .waitrequest
		.clock_cross_dma_to_pcie_s0_address                           (mm_interconnect_3_clock_cross_dma_to_pcie_s0_address),             //                             clock_cross_dma_to_pcie_s0.address
		.clock_cross_dma_to_pcie_s0_write                             (mm_interconnect_3_clock_cross_dma_to_pcie_s0_write),               //                                                       .write
		.clock_cross_dma_to_pcie_s0_read                              (mm_interconnect_3_clock_cross_dma_to_pcie_s0_read),                //                                                       .read
		.clock_cross_dma_to_pcie_s0_readdata                          (mm_interconnect_3_clock_cross_dma_to_pcie_s0_readdata),            //                                                       .readdata
		.clock_cross_dma_to_pcie_s0_writedata                         (mm_interconnect_3_clock_cross_dma_to_pcie_s0_writedata),           //                                                       .writedata
		.clock_cross_dma_to_pcie_s0_burstcount                        (mm_interconnect_3_clock_cross_dma_to_pcie_s0_burstcount),          //                                                       .burstcount
		.clock_cross_dma_to_pcie_s0_byteenable                        (mm_interconnect_3_clock_cross_dma_to_pcie_s0_byteenable),          //                                                       .byteenable
		.clock_cross_dma_to_pcie_s0_readdatavalid                     (mm_interconnect_3_clock_cross_dma_to_pcie_s0_readdatavalid),       //                                                       .readdatavalid
		.clock_cross_dma_to_pcie_s0_waitrequest                       (mm_interconnect_3_clock_cross_dma_to_pcie_s0_waitrequest),         //                                                       .waitrequest
		.clock_cross_dma_to_pcie_s0_debugaccess                       (mm_interconnect_3_clock_cross_dma_to_pcie_s0_debugaccess)          //                                                       .debugaccess
	);

	system_acl_iface_mm_interconnect_5 mm_interconnect_5 (
		.ddr3a_afi_clk_clk                                             (ddr3a_afi_clk_clk),                                   //                                           ddr3a_afi_clk.clk
		.clock_cross_kernel_mem_0_m0_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                  // clock_cross_kernel_mem_0_m0_reset_reset_bridge_in_reset.reset
		.em_pc_0_avl_in_translator_reset_reset_bridge_in_reset_reset   (reset_controller_ddr3a_reset_out_reset),              //   em_pc_0_avl_in_translator_reset_reset_bridge_in_reset.reset
		.em_pc_0_avl_reset_n_reset_bridge_in_reset_reset               (reset_controller_ddr3a_reset_out_reset),              //               em_pc_0_avl_reset_n_reset_bridge_in_reset.reset
		.clock_cross_kernel_mem_0_m0_address                           (clock_cross_kernel_mem_0_m0_address),                 //                             clock_cross_kernel_mem_0_m0.address
		.clock_cross_kernel_mem_0_m0_waitrequest                       (clock_cross_kernel_mem_0_m0_waitrequest),             //                                                        .waitrequest
		.clock_cross_kernel_mem_0_m0_burstcount                        (clock_cross_kernel_mem_0_m0_burstcount),              //                                                        .burstcount
		.clock_cross_kernel_mem_0_m0_byteenable                        (clock_cross_kernel_mem_0_m0_byteenable),              //                                                        .byteenable
		.clock_cross_kernel_mem_0_m0_read                              (clock_cross_kernel_mem_0_m0_read),                    //                                                        .read
		.clock_cross_kernel_mem_0_m0_readdata                          (clock_cross_kernel_mem_0_m0_readdata),                //                                                        .readdata
		.clock_cross_kernel_mem_0_m0_readdatavalid                     (clock_cross_kernel_mem_0_m0_readdatavalid),           //                                                        .readdatavalid
		.clock_cross_kernel_mem_0_m0_write                             (clock_cross_kernel_mem_0_m0_write),                   //                                                        .write
		.clock_cross_kernel_mem_0_m0_writedata                         (clock_cross_kernel_mem_0_m0_writedata),               //                                                        .writedata
		.clock_cross_kernel_mem_0_m0_debugaccess                       (clock_cross_kernel_mem_0_m0_debugaccess),             //                                                        .debugaccess
		.em_pc_0_avl_in_address                                        (mm_interconnect_5_em_pc_0_avl_in_address),            //                                          em_pc_0_avl_in.address
		.em_pc_0_avl_in_write                                          (mm_interconnect_5_em_pc_0_avl_in_write),              //                                                        .write
		.em_pc_0_avl_in_read                                           (mm_interconnect_5_em_pc_0_avl_in_read),               //                                                        .read
		.em_pc_0_avl_in_readdata                                       (mm_interconnect_5_em_pc_0_avl_in_readdata),           //                                                        .readdata
		.em_pc_0_avl_in_writedata                                      (mm_interconnect_5_em_pc_0_avl_in_writedata),          //                                                        .writedata
		.em_pc_0_avl_in_beginbursttransfer                             (mm_interconnect_5_em_pc_0_avl_in_beginbursttransfer), //                                                        .beginbursttransfer
		.em_pc_0_avl_in_burstcount                                     (mm_interconnect_5_em_pc_0_avl_in_burstcount),         //                                                        .burstcount
		.em_pc_0_avl_in_byteenable                                     (mm_interconnect_5_em_pc_0_avl_in_byteenable),         //                                                        .byteenable
		.em_pc_0_avl_in_readdatavalid                                  (mm_interconnect_5_em_pc_0_avl_in_readdatavalid),      //                                                        .readdatavalid
		.em_pc_0_avl_in_waitrequest                                    (mm_interconnect_5_em_pc_0_avl_in_waitrequest)         //                                                        .waitrequest
	);

	system_acl_iface_mm_interconnect_6 mm_interconnect_6 (
		.ddr3a_afi_clk_clk                                           (ddr3a_afi_clk_clk),                                         //                                         ddr3a_afi_clk.clk
		.acl_memory_bank_divider_0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                        // acl_memory_bank_divider_0_reset_reset_bridge_in_reset.reset
		.em_pc_0_avl_reset_n_reset_bridge_in_reset_reset             (reset_controller_ddr3a_reset_out_reset),                    //             em_pc_0_avl_reset_n_reset_bridge_in_reset.reset
		.pipe_stage_ddr3a_iface_reset_reset_bridge_in_reset_reset    (reset_controller_ddr3a_reset_out_reset),                    //    pipe_stage_ddr3a_iface_reset_reset_bridge_in_reset.reset
		.acl_memory_bank_divider_0_bank1_address                     (acl_memory_bank_divider_0_bank1_address),                   //                       acl_memory_bank_divider_0_bank1.address
		.acl_memory_bank_divider_0_bank1_waitrequest                 (acl_memory_bank_divider_0_bank1_waitrequest),               //                                                      .waitrequest
		.acl_memory_bank_divider_0_bank1_burstcount                  (acl_memory_bank_divider_0_bank1_burstcount),                //                                                      .burstcount
		.acl_memory_bank_divider_0_bank1_byteenable                  (acl_memory_bank_divider_0_bank1_byteenable),                //                                                      .byteenable
		.acl_memory_bank_divider_0_bank1_read                        (acl_memory_bank_divider_0_bank1_read),                      //                                                      .read
		.acl_memory_bank_divider_0_bank1_readdata                    (acl_memory_bank_divider_0_bank1_readdata),                  //                                                      .readdata
		.acl_memory_bank_divider_0_bank1_readdatavalid               (acl_memory_bank_divider_0_bank1_readdatavalid),             //                                                      .readdatavalid
		.acl_memory_bank_divider_0_bank1_write                       (acl_memory_bank_divider_0_bank1_write),                     //                                                      .write
		.acl_memory_bank_divider_0_bank1_writedata                   (acl_memory_bank_divider_0_bank1_writedata),                 //                                                      .writedata
		.em_pc_0_avl_out_address                                     (em_pc_0_avl_out_address),                                   //                                       em_pc_0_avl_out.address
		.em_pc_0_avl_out_waitrequest                                 (em_pc_0_avl_out_waitrequest),                               //                                                      .waitrequest
		.em_pc_0_avl_out_burstcount                                  (em_pc_0_avl_out_burstcount),                                //                                                      .burstcount
		.em_pc_0_avl_out_byteenable                                  (em_pc_0_avl_out_byteenable),                                //                                                      .byteenable
		.em_pc_0_avl_out_beginbursttransfer                          (em_pc_0_avl_out_beginbursttransfer),                        //                                                      .beginbursttransfer
		.em_pc_0_avl_out_read                                        (em_pc_0_avl_out_read),                                      //                                                      .read
		.em_pc_0_avl_out_readdata                                    (em_pc_0_avl_out_readdata),                                  //                                                      .readdata
		.em_pc_0_avl_out_readdatavalid                               (em_pc_0_avl_out_readdatavalid),                             //                                                      .readdatavalid
		.em_pc_0_avl_out_write                                       (em_pc_0_avl_out_write),                                     //                                                      .write
		.em_pc_0_avl_out_writedata                                   (em_pc_0_avl_out_writedata),                                 //                                                      .writedata
		.pipe_stage_ddr3a_iface_s0_address                           (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_address),       //                             pipe_stage_ddr3a_iface_s0.address
		.pipe_stage_ddr3a_iface_s0_write                             (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_write),         //                                                      .write
		.pipe_stage_ddr3a_iface_s0_read                              (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_read),          //                                                      .read
		.pipe_stage_ddr3a_iface_s0_readdata                          (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_readdata),      //                                                      .readdata
		.pipe_stage_ddr3a_iface_s0_writedata                         (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_writedata),     //                                                      .writedata
		.pipe_stage_ddr3a_iface_s0_burstcount                        (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_burstcount),    //                                                      .burstcount
		.pipe_stage_ddr3a_iface_s0_byteenable                        (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_byteenable),    //                                                      .byteenable
		.pipe_stage_ddr3a_iface_s0_readdatavalid                     (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_readdatavalid), //                                                      .readdatavalid
		.pipe_stage_ddr3a_iface_s0_waitrequest                       (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_waitrequest),   //                                                      .waitrequest
		.pipe_stage_ddr3a_iface_s0_debugaccess                       (mm_interconnect_6_pipe_stage_ddr3a_iface_s0_debugaccess)    //                                                      .debugaccess
	);

	system_acl_iface_mm_interconnect_7 mm_interconnect_7 (
		.ddr3b_afi_clk_clk                                             (ddr3b_afi_clk_clk),                                   //                                           ddr3b_afi_clk.clk
		.clock_cross_kernel_mem_1_m0_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                  // clock_cross_kernel_mem_1_m0_reset_reset_bridge_in_reset.reset
		.em_pc_1_avl_in_translator_reset_reset_bridge_in_reset_reset   (reset_controller_ddr3b_reset_out_reset),              //   em_pc_1_avl_in_translator_reset_reset_bridge_in_reset.reset
		.em_pc_1_avl_reset_n_reset_bridge_in_reset_reset               (reset_controller_ddr3b_reset_out_reset),              //               em_pc_1_avl_reset_n_reset_bridge_in_reset.reset
		.clock_cross_kernel_mem_1_m0_address                           (clock_cross_kernel_mem_1_m0_address),                 //                             clock_cross_kernel_mem_1_m0.address
		.clock_cross_kernel_mem_1_m0_waitrequest                       (clock_cross_kernel_mem_1_m0_waitrequest),             //                                                        .waitrequest
		.clock_cross_kernel_mem_1_m0_burstcount                        (clock_cross_kernel_mem_1_m0_burstcount),              //                                                        .burstcount
		.clock_cross_kernel_mem_1_m0_byteenable                        (clock_cross_kernel_mem_1_m0_byteenable),              //                                                        .byteenable
		.clock_cross_kernel_mem_1_m0_read                              (clock_cross_kernel_mem_1_m0_read),                    //                                                        .read
		.clock_cross_kernel_mem_1_m0_readdata                          (clock_cross_kernel_mem_1_m0_readdata),                //                                                        .readdata
		.clock_cross_kernel_mem_1_m0_readdatavalid                     (clock_cross_kernel_mem_1_m0_readdatavalid),           //                                                        .readdatavalid
		.clock_cross_kernel_mem_1_m0_write                             (clock_cross_kernel_mem_1_m0_write),                   //                                                        .write
		.clock_cross_kernel_mem_1_m0_writedata                         (clock_cross_kernel_mem_1_m0_writedata),               //                                                        .writedata
		.clock_cross_kernel_mem_1_m0_debugaccess                       (clock_cross_kernel_mem_1_m0_debugaccess),             //                                                        .debugaccess
		.em_pc_1_avl_in_address                                        (mm_interconnect_7_em_pc_1_avl_in_address),            //                                          em_pc_1_avl_in.address
		.em_pc_1_avl_in_write                                          (mm_interconnect_7_em_pc_1_avl_in_write),              //                                                        .write
		.em_pc_1_avl_in_read                                           (mm_interconnect_7_em_pc_1_avl_in_read),               //                                                        .read
		.em_pc_1_avl_in_readdata                                       (mm_interconnect_7_em_pc_1_avl_in_readdata),           //                                                        .readdata
		.em_pc_1_avl_in_writedata                                      (mm_interconnect_7_em_pc_1_avl_in_writedata),          //                                                        .writedata
		.em_pc_1_avl_in_beginbursttransfer                             (mm_interconnect_7_em_pc_1_avl_in_beginbursttransfer), //                                                        .beginbursttransfer
		.em_pc_1_avl_in_burstcount                                     (mm_interconnect_7_em_pc_1_avl_in_burstcount),         //                                                        .burstcount
		.em_pc_1_avl_in_byteenable                                     (mm_interconnect_7_em_pc_1_avl_in_byteenable),         //                                                        .byteenable
		.em_pc_1_avl_in_readdatavalid                                  (mm_interconnect_7_em_pc_1_avl_in_readdatavalid),      //                                                        .readdatavalid
		.em_pc_1_avl_in_waitrequest                                    (mm_interconnect_7_em_pc_1_avl_in_waitrequest)         //                                                        .waitrequest
	);

	system_acl_iface_mm_interconnect_8 mm_interconnect_8 (
		.pcie_coreclkout_clk                                        (pcie_coreclkout_clk),                                     //                                      pcie_coreclkout.clk
		.pcie_Rxm_BAR0_translator_reset_reset_bridge_in_reset_reset (rst_controller_008_reset_out_reset),                      // pcie_Rxm_BAR0_translator_reset_reset_bridge_in_reset.reset
		.pipe_stage_host_ctrl_reset_reset_bridge_in_reset_reset     (reset_controller_pcie_reset_out_reset),                   //     pipe_stage_host_ctrl_reset_reset_bridge_in_reset.reset
		.pcie_Rxm_BAR0_address                                      (pcie_rxm_bar0_address),                                   //                                        pcie_Rxm_BAR0.address
		.pcie_Rxm_BAR0_waitrequest                                  (pcie_rxm_bar0_waitrequest),                               //                                                     .waitrequest
		.pcie_Rxm_BAR0_burstcount                                   (pcie_rxm_bar0_burstcount),                                //                                                     .burstcount
		.pcie_Rxm_BAR0_byteenable                                   (pcie_rxm_bar0_byteenable),                                //                                                     .byteenable
		.pcie_Rxm_BAR0_read                                         (pcie_rxm_bar0_read),                                      //                                                     .read
		.pcie_Rxm_BAR0_readdata                                     (pcie_rxm_bar0_readdata),                                  //                                                     .readdata
		.pcie_Rxm_BAR0_readdatavalid                                (pcie_rxm_bar0_readdatavalid),                             //                                                     .readdatavalid
		.pcie_Rxm_BAR0_write                                        (pcie_rxm_bar0_write),                                     //                                                     .write
		.pcie_Rxm_BAR0_writedata                                    (pcie_rxm_bar0_writedata),                                 //                                                     .writedata
		.pipe_stage_host_ctrl_s0_address                            (mm_interconnect_8_pipe_stage_host_ctrl_s0_address),       //                              pipe_stage_host_ctrl_s0.address
		.pipe_stage_host_ctrl_s0_write                              (mm_interconnect_8_pipe_stage_host_ctrl_s0_write),         //                                                     .write
		.pipe_stage_host_ctrl_s0_read                               (mm_interconnect_8_pipe_stage_host_ctrl_s0_read),          //                                                     .read
		.pipe_stage_host_ctrl_s0_readdata                           (mm_interconnect_8_pipe_stage_host_ctrl_s0_readdata),      //                                                     .readdata
		.pipe_stage_host_ctrl_s0_writedata                          (mm_interconnect_8_pipe_stage_host_ctrl_s0_writedata),     //                                                     .writedata
		.pipe_stage_host_ctrl_s0_burstcount                         (mm_interconnect_8_pipe_stage_host_ctrl_s0_burstcount),    //                                                     .burstcount
		.pipe_stage_host_ctrl_s0_byteenable                         (mm_interconnect_8_pipe_stage_host_ctrl_s0_byteenable),    //                                                     .byteenable
		.pipe_stage_host_ctrl_s0_readdatavalid                      (mm_interconnect_8_pipe_stage_host_ctrl_s0_readdatavalid), //                                                     .readdatavalid
		.pipe_stage_host_ctrl_s0_waitrequest                        (mm_interconnect_8_pipe_stage_host_ctrl_s0_waitrequest),   //                                                     .waitrequest
		.pipe_stage_host_ctrl_s0_debugaccess                        (mm_interconnect_8_pipe_stage_host_ctrl_s0_debugaccess)    //                                                     .debugaccess
	);

	system_acl_iface_mm_interconnect_9 mm_interconnect_9 (
		.pcie_coreclkout_clk                                          (pcie_coreclkout_clk),                      //                                        pcie_coreclkout.clk
		.clock_cross_dma_to_pcie_m0_reset_reset_bridge_in_reset_reset (reset_controller_pcie_reset_out_reset),    // clock_cross_dma_to_pcie_m0_reset_reset_bridge_in_reset.reset
		.pcie_Txs_translator_reset_reset_bridge_in_reset_reset        (rst_controller_008_reset_out_reset),       //        pcie_Txs_translator_reset_reset_bridge_in_reset.reset
		.clock_cross_dma_to_pcie_m0_address                           (clock_cross_dma_to_pcie_m0_address),       //                             clock_cross_dma_to_pcie_m0.address
		.clock_cross_dma_to_pcie_m0_waitrequest                       (clock_cross_dma_to_pcie_m0_waitrequest),   //                                                       .waitrequest
		.clock_cross_dma_to_pcie_m0_burstcount                        (clock_cross_dma_to_pcie_m0_burstcount),    //                                                       .burstcount
		.clock_cross_dma_to_pcie_m0_byteenable                        (clock_cross_dma_to_pcie_m0_byteenable),    //                                                       .byteenable
		.clock_cross_dma_to_pcie_m0_read                              (clock_cross_dma_to_pcie_m0_read),          //                                                       .read
		.clock_cross_dma_to_pcie_m0_readdata                          (clock_cross_dma_to_pcie_m0_readdata),      //                                                       .readdata
		.clock_cross_dma_to_pcie_m0_readdatavalid                     (clock_cross_dma_to_pcie_m0_readdatavalid), //                                                       .readdatavalid
		.clock_cross_dma_to_pcie_m0_write                             (clock_cross_dma_to_pcie_m0_write),         //                                                       .write
		.clock_cross_dma_to_pcie_m0_writedata                         (clock_cross_dma_to_pcie_m0_writedata),     //                                                       .writedata
		.clock_cross_dma_to_pcie_m0_debugaccess                       (clock_cross_dma_to_pcie_m0_debugaccess),   //                                                       .debugaccess
		.pcie_Txs_address                                             (mm_interconnect_9_pcie_txs_address),       //                                               pcie_Txs.address
		.pcie_Txs_write                                               (mm_interconnect_9_pcie_txs_write),         //                                                       .write
		.pcie_Txs_read                                                (mm_interconnect_9_pcie_txs_read),          //                                                       .read
		.pcie_Txs_readdata                                            (mm_interconnect_9_pcie_txs_readdata),      //                                                       .readdata
		.pcie_Txs_writedata                                           (mm_interconnect_9_pcie_txs_writedata),     //                                                       .writedata
		.pcie_Txs_burstcount                                          (mm_interconnect_9_pcie_txs_burstcount),    //                                                       .burstcount
		.pcie_Txs_byteenable                                          (mm_interconnect_9_pcie_txs_byteenable),    //                                                       .byteenable
		.pcie_Txs_readdatavalid                                       (mm_interconnect_9_pcie_txs_readdatavalid), //                                                       .readdatavalid
		.pcie_Txs_waitrequest                                         (mm_interconnect_9_pcie_txs_waitrequest),   //                                                       .waitrequest
		.pcie_Txs_chipselect                                          (mm_interconnect_9_pcie_txs_chipselect)     //                                                       .chipselect
	);

	system_acl_iface_mm_interconnect_10 mm_interconnect_10 (
		.ddr3b_afi_clk_clk                                             (ddr3b_afi_clk_clk),                                          //                                           ddr3b_afi_clk.clk
		.clock_cross_dma_to_ddr3b_m0_reset_reset_bridge_in_reset_reset (reset_controller_ddr3b_reset_out_reset),                     // clock_cross_dma_to_ddr3b_m0_reset_reset_bridge_in_reset.reset
		.em_pc_1_avl_reset_n_reset_bridge_in_reset_reset               (reset_controller_ddr3b_reset_out_reset),                     //               em_pc_1_avl_reset_n_reset_bridge_in_reset.reset
		.clock_cross_dma_to_ddr3b_m0_address                           (clock_cross_dma_to_ddr3b_m0_address),                        //                             clock_cross_dma_to_ddr3b_m0.address
		.clock_cross_dma_to_ddr3b_m0_waitrequest                       (clock_cross_dma_to_ddr3b_m0_waitrequest),                    //                                                        .waitrequest
		.clock_cross_dma_to_ddr3b_m0_burstcount                        (clock_cross_dma_to_ddr3b_m0_burstcount),                     //                                                        .burstcount
		.clock_cross_dma_to_ddr3b_m0_byteenable                        (clock_cross_dma_to_ddr3b_m0_byteenable),                     //                                                        .byteenable
		.clock_cross_dma_to_ddr3b_m0_read                              (clock_cross_dma_to_ddr3b_m0_read),                           //                                                        .read
		.clock_cross_dma_to_ddr3b_m0_readdata                          (clock_cross_dma_to_ddr3b_m0_readdata),                       //                                                        .readdata
		.clock_cross_dma_to_ddr3b_m0_readdatavalid                     (clock_cross_dma_to_ddr3b_m0_readdatavalid),                  //                                                        .readdatavalid
		.clock_cross_dma_to_ddr3b_m0_write                             (clock_cross_dma_to_ddr3b_m0_write),                          //                                                        .write
		.clock_cross_dma_to_ddr3b_m0_writedata                         (clock_cross_dma_to_ddr3b_m0_writedata),                      //                                                        .writedata
		.clock_cross_dma_to_ddr3b_m0_debugaccess                       (clock_cross_dma_to_ddr3b_m0_debugaccess),                    //                                                        .debugaccess
		.em_pc_1_avl_out_address                                       (em_pc_1_avl_out_address),                                    //                                         em_pc_1_avl_out.address
		.em_pc_1_avl_out_waitrequest                                   (em_pc_1_avl_out_waitrequest),                                //                                                        .waitrequest
		.em_pc_1_avl_out_burstcount                                    (em_pc_1_avl_out_burstcount),                                 //                                                        .burstcount
		.em_pc_1_avl_out_byteenable                                    (em_pc_1_avl_out_byteenable),                                 //                                                        .byteenable
		.em_pc_1_avl_out_beginbursttransfer                            (em_pc_1_avl_out_beginbursttransfer),                         //                                                        .beginbursttransfer
		.em_pc_1_avl_out_read                                          (em_pc_1_avl_out_read),                                       //                                                        .read
		.em_pc_1_avl_out_readdata                                      (em_pc_1_avl_out_readdata),                                   //                                                        .readdata
		.em_pc_1_avl_out_readdatavalid                                 (em_pc_1_avl_out_readdatavalid),                              //                                                        .readdatavalid
		.em_pc_1_avl_out_write                                         (em_pc_1_avl_out_write),                                      //                                                        .write
		.em_pc_1_avl_out_writedata                                     (em_pc_1_avl_out_writedata),                                  //                                                        .writedata
		.pipe_stage_ddr3b_iface_s0_address                             (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_address),       //                               pipe_stage_ddr3b_iface_s0.address
		.pipe_stage_ddr3b_iface_s0_write                               (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_write),         //                                                        .write
		.pipe_stage_ddr3b_iface_s0_read                                (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_read),          //                                                        .read
		.pipe_stage_ddr3b_iface_s0_readdata                            (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_readdata),      //                                                        .readdata
		.pipe_stage_ddr3b_iface_s0_writedata                           (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_writedata),     //                                                        .writedata
		.pipe_stage_ddr3b_iface_s0_burstcount                          (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_burstcount),    //                                                        .burstcount
		.pipe_stage_ddr3b_iface_s0_byteenable                          (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_byteenable),    //                                                        .byteenable
		.pipe_stage_ddr3b_iface_s0_readdatavalid                       (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_readdatavalid), //                                                        .readdatavalid
		.pipe_stage_ddr3b_iface_s0_waitrequest                         (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_waitrequest),   //                                                        .waitrequest
		.pipe_stage_ddr3b_iface_s0_debugaccess                         (mm_interconnect_10_pipe_stage_ddr3b_iface_s0_debugaccess)    //                                                        .debugaccess
	);

	system_acl_iface_mm_interconnect_12 mm_interconnect_12 (
		.ddr3a_afi_clk_clk                                             (ddr3a_afi_clk_clk),                                            //                                           ddr3a_afi_clk.clk
		.acl_memory_bank_divider_0_reset_reset_bridge_in_reset_reset   (rst_controller_002_reset_out_reset),                           //   acl_memory_bank_divider_0_reset_reset_bridge_in_reset.reset
		.clock_cross_dma_to_ddr3b_s0_reset_reset_bridge_in_reset_reset (reset_controller_ddr3a_reset_out_reset),                       // clock_cross_dma_to_ddr3b_s0_reset_reset_bridge_in_reset.reset
		.acl_memory_bank_divider_0_bank2_address                       (acl_memory_bank_divider_0_bank2_address),                      //                         acl_memory_bank_divider_0_bank2.address
		.acl_memory_bank_divider_0_bank2_waitrequest                   (acl_memory_bank_divider_0_bank2_waitrequest),                  //                                                        .waitrequest
		.acl_memory_bank_divider_0_bank2_burstcount                    (acl_memory_bank_divider_0_bank2_burstcount),                   //                                                        .burstcount
		.acl_memory_bank_divider_0_bank2_byteenable                    (acl_memory_bank_divider_0_bank2_byteenable),                   //                                                        .byteenable
		.acl_memory_bank_divider_0_bank2_read                          (acl_memory_bank_divider_0_bank2_read),                         //                                                        .read
		.acl_memory_bank_divider_0_bank2_readdata                      (acl_memory_bank_divider_0_bank2_readdata),                     //                                                        .readdata
		.acl_memory_bank_divider_0_bank2_readdatavalid                 (acl_memory_bank_divider_0_bank2_readdatavalid),                //                                                        .readdatavalid
		.acl_memory_bank_divider_0_bank2_write                         (acl_memory_bank_divider_0_bank2_write),                        //                                                        .write
		.acl_memory_bank_divider_0_bank2_writedata                     (acl_memory_bank_divider_0_bank2_writedata),                    //                                                        .writedata
		.clock_cross_dma_to_ddr3b_s0_address                           (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_address),       //                             clock_cross_dma_to_ddr3b_s0.address
		.clock_cross_dma_to_ddr3b_s0_write                             (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_write),         //                                                        .write
		.clock_cross_dma_to_ddr3b_s0_read                              (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_read),          //                                                        .read
		.clock_cross_dma_to_ddr3b_s0_readdata                          (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_readdata),      //                                                        .readdata
		.clock_cross_dma_to_ddr3b_s0_writedata                         (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_writedata),     //                                                        .writedata
		.clock_cross_dma_to_ddr3b_s0_burstcount                        (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_burstcount),    //                                                        .burstcount
		.clock_cross_dma_to_ddr3b_s0_byteenable                        (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_byteenable),    //                                                        .byteenable
		.clock_cross_dma_to_ddr3b_s0_readdatavalid                     (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_readdatavalid), //                                                        .readdatavalid
		.clock_cross_dma_to_ddr3b_s0_waitrequest                       (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_waitrequest),   //                                                        .waitrequest
		.clock_cross_dma_to_ddr3b_s0_debugaccess                       (mm_interconnect_12_clock_cross_dma_to_ddr3b_s0_debugaccess)    //                                                        .debugaccess
	);

	system_acl_iface_irq_mapper irq_mapper (
		.clk           (pcie_coreclkout_clk),                //       clk.clk
		.reset         (rst_controller_008_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (pcie_rxmirq_irq)                     //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (kernel_clk_clk),                     //       receiver_clk.clk
		.sender_clk     (pcie_coreclkout_clk),                //         sender_clk.clk
		.receiver_reset (rst_controller_009_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_008_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (ddr3a_afi_clk_clk),                  //       receiver_clk.clk
		.sender_clk     (pcie_coreclkout_clk),                //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_008_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_controller_global_reset_out_reset), // reset_in0.reset
		.clk            (ddr3a_afi_clk_clk),                       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),          // reset_out.reset
		.reset_req      (),                                        // (terminated)
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_in1      (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (reset_controller_global_reset_out_reset), // reset_in0.reset
		.clk            (temperature_pll_outclk0_clk),             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),      // reset_out.reset
		.reset_req      (),                                        // (terminated)
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_in1      (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (reset_controller_ddr3b_reset_out_reset), // reset_in0.reset
		.clk            (ddr3a_afi_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~kernel_interface_sw_reset_export_reset), // reset_in0.reset
		.clk            (ddr3a_afi_clk_clk),                       //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),      // reset_out.reset
		.reset_req      (),                                        // (terminated)
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_in1      (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~kernel_interface_sw_reset_export_reset), // reset_in0.reset
		.clk            (ddr3b_afi_clk_clk),                       //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),      // reset_out.reset
		.reset_req      (),                                        // (terminated)
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_in1      (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_n),                           // reset_in0.reset
		.clk            (config_clk_clk),                     //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (reset_controller_global_reset_out_reset), // reset_in0.reset
		.clk            (pcie_coreclkout_clk),                     //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset),      // reset_out.reset
		.reset_req      (),                                        // (terminated)
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_in1      (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (reset_controller_global_reset_out_reset), // reset_in0.reset
		.clk            (ddr3b_afi_clk_clk),                       //       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset),      // reset_out.reset
		.reset_req      (),                                        // (terminated)
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_in1      (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_008 (
		.reset_in0      (~pcie_nreset_status_reset),          // reset_in0.reset
		.clk            (pcie_coreclkout_clk),                //       clk.clk
		.reset_out      (rst_controller_008_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_009 (
		.reset_in0      (reset_controller_pcie_reset_out_reset), // reset_in0.reset
		.clk            (kernel_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_009_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                      // (terminated)
		.reset_req_in0  (1'b0),                                  // (terminated)
		.reset_in1      (1'b0),                                  // (terminated)
		.reset_req_in1  (1'b0),                                  // (terminated)
		.reset_in2      (1'b0),                                  // (terminated)
		.reset_req_in2  (1'b0),                                  // (terminated)
		.reset_in3      (1'b0),                                  // (terminated)
		.reset_req_in3  (1'b0),                                  // (terminated)
		.reset_in4      (1'b0),                                  // (terminated)
		.reset_req_in4  (1'b0),                                  // (terminated)
		.reset_in5      (1'b0),                                  // (terminated)
		.reset_req_in5  (1'b0),                                  // (terminated)
		.reset_in6      (1'b0),                                  // (terminated)
		.reset_req_in6  (1'b0),                                  // (terminated)
		.reset_in7      (1'b0),                                  // (terminated)
		.reset_req_in7  (1'b0),                                  // (terminated)
		.reset_in8      (1'b0),                                  // (terminated)
		.reset_req_in8  (1'b0),                                  // (terminated)
		.reset_in9      (1'b0),                                  // (terminated)
		.reset_req_in9  (1'b0),                                  // (terminated)
		.reset_in10     (1'b0),                                  // (terminated)
		.reset_req_in10 (1'b0),                                  // (terminated)
		.reset_in11     (1'b0),                                  // (terminated)
		.reset_req_in11 (1'b0),                                  // (terminated)
		.reset_in12     (1'b0),                                  // (terminated)
		.reset_req_in12 (1'b0),                                  // (terminated)
		.reset_in13     (1'b0),                                  // (terminated)
		.reset_req_in13 (1'b0),                                  // (terminated)
		.reset_in14     (1'b0),                                  // (terminated)
		.reset_req_in14 (1'b0),                                  // (terminated)
		.reset_in15     (1'b0),                                  // (terminated)
		.reset_req_in15 (1'b0)                                   // (terminated)
	);

endmodule

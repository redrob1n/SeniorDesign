// system.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module system (
		input  wire         config_clk_clk,                        //         config_clk.clk
		output wire [14:0]  ddr3a_mem_a,                           //              ddr3a.mem_a
		output wire [2:0]   ddr3a_mem_ba,                          //                   .mem_ba
		output wire [0:0]   ddr3a_mem_ck,                          //                   .mem_ck
		output wire [0:0]   ddr3a_mem_ck_n,                        //                   .mem_ck_n
		output wire [0:0]   ddr3a_mem_cke,                         //                   .mem_cke
		output wire [0:0]   ddr3a_mem_cs_n,                        //                   .mem_cs_n
		output wire [7:0]   ddr3a_mem_dm,                          //                   .mem_dm
		output wire [0:0]   ddr3a_mem_ras_n,                       //                   .mem_ras_n
		output wire [0:0]   ddr3a_mem_cas_n,                       //                   .mem_cas_n
		output wire [0:0]   ddr3a_mem_we_n,                        //                   .mem_we_n
		output wire         ddr3a_mem_reset_n,                     //                   .mem_reset_n
		inout  wire [63:0]  ddr3a_mem_dq,                          //                   .mem_dq
		inout  wire [7:0]   ddr3a_mem_dqs,                         //                   .mem_dqs
		inout  wire [7:0]   ddr3a_mem_dqs_n,                       //                   .mem_dqs_n
		output wire [0:0]   ddr3a_mem_odt,                         //                   .mem_odt
		input  wire         ddr3a_mem_oct_rzqin,                   //      ddr3a_mem_oct.rzqin
		input  wire         ddr3a_pll_ref_clk,                     //      ddr3a_pll_ref.clk
		output wire [14:0]  ddr3b_mem_a,                           //              ddr3b.mem_a
		output wire [2:0]   ddr3b_mem_ba,                          //                   .mem_ba
		output wire [0:0]   ddr3b_mem_ck,                          //                   .mem_ck
		output wire [0:0]   ddr3b_mem_ck_n,                        //                   .mem_ck_n
		output wire [0:0]   ddr3b_mem_cke,                         //                   .mem_cke
		output wire [0:0]   ddr3b_mem_cs_n,                        //                   .mem_cs_n
		output wire [7:0]   ddr3b_mem_dm,                          //                   .mem_dm
		output wire [0:0]   ddr3b_mem_ras_n,                       //                   .mem_ras_n
		output wire [0:0]   ddr3b_mem_cas_n,                       //                   .mem_cas_n
		output wire [0:0]   ddr3b_mem_we_n,                        //                   .mem_we_n
		output wire         ddr3b_mem_reset_n,                     //                   .mem_reset_n
		inout  wire [63:0]  ddr3b_mem_dq,                          //                   .mem_dq
		inout  wire [7:0]   ddr3b_mem_dqs,                         //                   .mem_dqs
		inout  wire [7:0]   ddr3b_mem_dqs_n,                       //                   .mem_dqs_n
		output wire [0:0]   ddr3b_mem_odt,                         //                   .mem_odt
		input  wire         ddr3b_mem_oct_rzqin,                   //      ddr3b_mem_oct.rzqin
		input  wire         ddr3b_pll_ref_clk,                     //      ddr3b_pll_ref.clk
		input  wire         global_reset_reset_n,                  //       global_reset.reset_n
		input  wire         kernel_pll_refclk_clk,                 //  kernel_pll_refclk.clk
		input  wire         pcie_rx_in0,                           //               pcie.rx_in0
		input  wire         pcie_rx_in1,                           //                   .rx_in1
		input  wire         pcie_rx_in2,                           //                   .rx_in2
		input  wire         pcie_rx_in3,                           //                   .rx_in3
		input  wire         pcie_rx_in4,                           //                   .rx_in4
		input  wire         pcie_rx_in5,                           //                   .rx_in5
		input  wire         pcie_rx_in6,                           //                   .rx_in6
		input  wire         pcie_rx_in7,                           //                   .rx_in7
		output wire         pcie_tx_out0,                          //                   .tx_out0
		output wire         pcie_tx_out1,                          //                   .tx_out1
		output wire         pcie_tx_out2,                          //                   .tx_out2
		output wire         pcie_tx_out3,                          //                   .tx_out3
		output wire         pcie_tx_out4,                          //                   .tx_out4
		output wire         pcie_tx_out5,                          //                   .tx_out5
		output wire         pcie_tx_out6,                          //                   .tx_out6
		output wire         pcie_tx_out7,                          //                   .tx_out7
		input  wire         pcie_npor_npor,                        //          pcie_npor.npor
		input  wire         pcie_npor_pin_perst,                   //                   .pin_perst
		output wire         pcie_npor_out_reset_n,                 //      pcie_npor_out.reset_n
		input  wire         pcie_refclk_clk,                       //        pcie_refclk.clk
		output wire [459:0] reconfig_from_xcvr_reconfig_from_xcvr, // reconfig_from_xcvr.reconfig_from_xcvr
		input  wire [699:0] reconfig_to_xcvr_reconfig_to_xcvr      //   reconfig_to_xcvr.reconfig_to_xcvr
	);

	wire   [63:0] avs_vadd_cra_cra_ring_cra_master_readdata;                       // genetic_algorithm_system:avs_vadd_cra_readdata -> avs_vadd_cra_cra_ring:avm_readdata
	wire          avs_vadd_cra_cra_ring_cra_master_read;                           // avs_vadd_cra_cra_ring:avm_read -> genetic_algorithm_system:avs_vadd_cra_read
	wire    [3:0] avs_vadd_cra_cra_ring_cra_master_address;                        // avs_vadd_cra_cra_ring:avm_addr -> genetic_algorithm_system:avs_vadd_cra_address
	wire    [7:0] avs_vadd_cra_cra_ring_cra_master_byteenable;                     // avs_vadd_cra_cra_ring:avm_byteena -> genetic_algorithm_system:avs_vadd_cra_byteenable
	wire          avs_vadd_cra_cra_ring_cra_master_readdatavalid;                  // genetic_algorithm_system:avs_vadd_cra_readdatavalid -> avs_vadd_cra_cra_ring:avm_readdatavalid
	wire          avs_vadd_cra_cra_ring_cra_master_write;                          // avs_vadd_cra_cra_ring:avm_write -> genetic_algorithm_system:avs_vadd_cra_write
	wire   [63:0] avs_vadd_cra_cra_ring_cra_master_writedata;                      // avs_vadd_cra_cra_ring:avm_writedata -> genetic_algorithm_system:avs_vadd_cra_writedata
	wire          acl_iface_kernel_clk_clk;                                        // acl_iface:kernel_clk_clk -> [avs_vadd_cra_cra_ring:clk, cra_root:clk, genetic_algorithm_system:clock, irq_mapper:clk, mm_interconnect_0:acl_iface_kernel_clk_clk, mm_interconnect_1:acl_iface_kernel_clk_clk, mm_interconnect_3:acl_iface_kernel_clk_clk, rst_controller:clk]
	wire          acl_iface_kernel_clk2x_clk;                                      // acl_iface:kernel_clk2x_clk -> genetic_algorithm_system:clock2x
	wire          cra_root_ring_out_datavalid;                                     // cra_root:ro_datavalid -> avs_vadd_cra_cra_ring:ri_datavalid
	wire          cra_root_ring_out_read;                                          // cra_root:ro_read -> avs_vadd_cra_cra_ring:ri_read
	wire   [63:0] cra_root_ring_out_data;                                          // cra_root:ro_data -> avs_vadd_cra_cra_ring:ri_data
	wire    [3:0] cra_root_ring_out_addr;                                          // cra_root:ro_addr -> avs_vadd_cra_cra_ring:ri_addr
	wire          cra_root_ring_out_write;                                         // cra_root:ro_write -> avs_vadd_cra_cra_ring:ri_write
	wire    [7:0] cra_root_ring_out_byteena;                                       // cra_root:ro_byteena -> avs_vadd_cra_cra_ring:ri_byteena
	wire          avs_vadd_cra_cra_ring_ring_out_datavalid;                        // avs_vadd_cra_cra_ring:ro_datavalid -> cra_root:ri_datavalid
	wire          avs_vadd_cra_cra_ring_ring_out_read;                             // avs_vadd_cra_cra_ring:ro_read -> cra_root:ri_read
	wire   [63:0] avs_vadd_cra_cra_ring_ring_out_data;                             // avs_vadd_cra_cra_ring:ro_data -> cra_root:ri_data
	wire    [3:0] avs_vadd_cra_cra_ring_ring_out_addr;                             // avs_vadd_cra_cra_ring:ro_addr -> cra_root:ri_addr
	wire          avs_vadd_cra_cra_ring_ring_out_write;                            // avs_vadd_cra_cra_ring:ro_write -> cra_root:ri_write
	wire    [7:0] avs_vadd_cra_cra_ring_ring_out_byteena;                          // avs_vadd_cra_cra_ring:ro_byteena -> cra_root:ri_byteena
	wire          acl_iface_kernel_reset_reset;                                    // acl_iface:kernel_reset_reset_n -> [avs_vadd_cra_cra_ring:rst_n, cra_root:rst_n, genetic_algorithm_system:resetn, mm_interconnect_0:genetic_algorithm_system_clock_reset_reset_reset_bridge_in_reset_reset, mm_interconnect_1:genetic_algorithm_system_clock_reset_reset_reset_bridge_in_reset_reset, mm_interconnect_3:cra_root_reset_reset_bridge_in_reset_reset]
	wire  [511:0] genetic_algorithm_system_avm_memgmem0_port_0_0_rw_readdata;      // mm_interconnect_0:genetic_algorithm_system_avm_memgmem0_port_0_0_rw_readdata -> genetic_algorithm_system:avm_memgmem0_port_0_0_rw_readdata
	wire          genetic_algorithm_system_avm_memgmem0_port_0_0_rw_waitrequest;   // mm_interconnect_0:genetic_algorithm_system_avm_memgmem0_port_0_0_rw_waitrequest -> genetic_algorithm_system:avm_memgmem0_port_0_0_rw_waitrequest
	wire   [30:0] genetic_algorithm_system_avm_memgmem0_port_0_0_rw_address;       // genetic_algorithm_system:avm_memgmem0_port_0_0_rw_address -> mm_interconnect_0:genetic_algorithm_system_avm_memgmem0_port_0_0_rw_address
	wire          genetic_algorithm_system_avm_memgmem0_port_0_0_rw_read;          // genetic_algorithm_system:avm_memgmem0_port_0_0_rw_read -> mm_interconnect_0:genetic_algorithm_system_avm_memgmem0_port_0_0_rw_read
	wire   [63:0] genetic_algorithm_system_avm_memgmem0_port_0_0_rw_byteenable;    // genetic_algorithm_system:avm_memgmem0_port_0_0_rw_byteenable -> mm_interconnect_0:genetic_algorithm_system_avm_memgmem0_port_0_0_rw_byteenable
	wire          genetic_algorithm_system_avm_memgmem0_port_0_0_rw_readdatavalid; // mm_interconnect_0:genetic_algorithm_system_avm_memgmem0_port_0_0_rw_readdatavalid -> genetic_algorithm_system:avm_memgmem0_port_0_0_rw_readdatavalid
	wire          genetic_algorithm_system_avm_memgmem0_port_0_0_rw_write;         // genetic_algorithm_system:avm_memgmem0_port_0_0_rw_write -> mm_interconnect_0:genetic_algorithm_system_avm_memgmem0_port_0_0_rw_write
	wire  [511:0] genetic_algorithm_system_avm_memgmem0_port_0_0_rw_writedata;     // genetic_algorithm_system:avm_memgmem0_port_0_0_rw_writedata -> mm_interconnect_0:genetic_algorithm_system_avm_memgmem0_port_0_0_rw_writedata
	wire    [4:0] genetic_algorithm_system_avm_memgmem0_port_0_0_rw_burstcount;    // genetic_algorithm_system:avm_memgmem0_port_0_0_rw_burstcount -> mm_interconnect_0:genetic_algorithm_system_avm_memgmem0_port_0_0_rw_burstcount
	wire  [511:0] mm_interconnect_0_acl_iface_kernel_mem0_readdata;                // acl_iface:kernel_mem0_readdata -> mm_interconnect_0:acl_iface_kernel_mem0_readdata
	wire          mm_interconnect_0_acl_iface_kernel_mem0_waitrequest;             // acl_iface:kernel_mem0_waitrequest -> mm_interconnect_0:acl_iface_kernel_mem0_waitrequest
	wire          mm_interconnect_0_acl_iface_kernel_mem0_debugaccess;             // mm_interconnect_0:acl_iface_kernel_mem0_debugaccess -> acl_iface:kernel_mem0_debugaccess
	wire   [30:0] mm_interconnect_0_acl_iface_kernel_mem0_address;                 // mm_interconnect_0:acl_iface_kernel_mem0_address -> acl_iface:kernel_mem0_address
	wire          mm_interconnect_0_acl_iface_kernel_mem0_read;                    // mm_interconnect_0:acl_iface_kernel_mem0_read -> acl_iface:kernel_mem0_read
	wire   [63:0] mm_interconnect_0_acl_iface_kernel_mem0_byteenable;              // mm_interconnect_0:acl_iface_kernel_mem0_byteenable -> acl_iface:kernel_mem0_byteenable
	wire          mm_interconnect_0_acl_iface_kernel_mem0_readdatavalid;           // acl_iface:kernel_mem0_readdatavalid -> mm_interconnect_0:acl_iface_kernel_mem0_readdatavalid
	wire          mm_interconnect_0_acl_iface_kernel_mem0_write;                   // mm_interconnect_0:acl_iface_kernel_mem0_write -> acl_iface:kernel_mem0_write
	wire  [511:0] mm_interconnect_0_acl_iface_kernel_mem0_writedata;               // mm_interconnect_0:acl_iface_kernel_mem0_writedata -> acl_iface:kernel_mem0_writedata
	wire    [4:0] mm_interconnect_0_acl_iface_kernel_mem0_burstcount;              // mm_interconnect_0:acl_iface_kernel_mem0_burstcount -> acl_iface:kernel_mem0_burstcount
	wire  [511:0] genetic_algorithm_system_avm_memgmem0_port_1_0_rw_readdata;      // mm_interconnect_1:genetic_algorithm_system_avm_memgmem0_port_1_0_rw_readdata -> genetic_algorithm_system:avm_memgmem0_port_1_0_rw_readdata
	wire          genetic_algorithm_system_avm_memgmem0_port_1_0_rw_waitrequest;   // mm_interconnect_1:genetic_algorithm_system_avm_memgmem0_port_1_0_rw_waitrequest -> genetic_algorithm_system:avm_memgmem0_port_1_0_rw_waitrequest
	wire   [30:0] genetic_algorithm_system_avm_memgmem0_port_1_0_rw_address;       // genetic_algorithm_system:avm_memgmem0_port_1_0_rw_address -> mm_interconnect_1:genetic_algorithm_system_avm_memgmem0_port_1_0_rw_address
	wire          genetic_algorithm_system_avm_memgmem0_port_1_0_rw_read;          // genetic_algorithm_system:avm_memgmem0_port_1_0_rw_read -> mm_interconnect_1:genetic_algorithm_system_avm_memgmem0_port_1_0_rw_read
	wire   [63:0] genetic_algorithm_system_avm_memgmem0_port_1_0_rw_byteenable;    // genetic_algorithm_system:avm_memgmem0_port_1_0_rw_byteenable -> mm_interconnect_1:genetic_algorithm_system_avm_memgmem0_port_1_0_rw_byteenable
	wire          genetic_algorithm_system_avm_memgmem0_port_1_0_rw_readdatavalid; // mm_interconnect_1:genetic_algorithm_system_avm_memgmem0_port_1_0_rw_readdatavalid -> genetic_algorithm_system:avm_memgmem0_port_1_0_rw_readdatavalid
	wire          genetic_algorithm_system_avm_memgmem0_port_1_0_rw_write;         // genetic_algorithm_system:avm_memgmem0_port_1_0_rw_write -> mm_interconnect_1:genetic_algorithm_system_avm_memgmem0_port_1_0_rw_write
	wire  [511:0] genetic_algorithm_system_avm_memgmem0_port_1_0_rw_writedata;     // genetic_algorithm_system:avm_memgmem0_port_1_0_rw_writedata -> mm_interconnect_1:genetic_algorithm_system_avm_memgmem0_port_1_0_rw_writedata
	wire    [4:0] genetic_algorithm_system_avm_memgmem0_port_1_0_rw_burstcount;    // genetic_algorithm_system:avm_memgmem0_port_1_0_rw_burstcount -> mm_interconnect_1:genetic_algorithm_system_avm_memgmem0_port_1_0_rw_burstcount
	wire  [511:0] mm_interconnect_1_acl_iface_kernel_mem1_readdata;                // acl_iface:kernel_mem1_readdata -> mm_interconnect_1:acl_iface_kernel_mem1_readdata
	wire          mm_interconnect_1_acl_iface_kernel_mem1_waitrequest;             // acl_iface:kernel_mem1_waitrequest -> mm_interconnect_1:acl_iface_kernel_mem1_waitrequest
	wire          mm_interconnect_1_acl_iface_kernel_mem1_debugaccess;             // mm_interconnect_1:acl_iface_kernel_mem1_debugaccess -> acl_iface:kernel_mem1_debugaccess
	wire   [30:0] mm_interconnect_1_acl_iface_kernel_mem1_address;                 // mm_interconnect_1:acl_iface_kernel_mem1_address -> acl_iface:kernel_mem1_address
	wire          mm_interconnect_1_acl_iface_kernel_mem1_read;                    // mm_interconnect_1:acl_iface_kernel_mem1_read -> acl_iface:kernel_mem1_read
	wire   [63:0] mm_interconnect_1_acl_iface_kernel_mem1_byteenable;              // mm_interconnect_1:acl_iface_kernel_mem1_byteenable -> acl_iface:kernel_mem1_byteenable
	wire          mm_interconnect_1_acl_iface_kernel_mem1_readdatavalid;           // acl_iface:kernel_mem1_readdatavalid -> mm_interconnect_1:acl_iface_kernel_mem1_readdatavalid
	wire          mm_interconnect_1_acl_iface_kernel_mem1_write;                   // mm_interconnect_1:acl_iface_kernel_mem1_write -> acl_iface:kernel_mem1_write
	wire  [511:0] mm_interconnect_1_acl_iface_kernel_mem1_writedata;               // mm_interconnect_1:acl_iface_kernel_mem1_writedata -> acl_iface:kernel_mem1_writedata
	wire    [4:0] mm_interconnect_1_acl_iface_kernel_mem1_burstcount;              // mm_interconnect_1:acl_iface_kernel_mem1_burstcount -> acl_iface:kernel_mem1_burstcount
	wire          acl_iface_kernel_cra_waitrequest;                                // mm_interconnect_3:acl_iface_kernel_cra_waitrequest -> acl_iface:kernel_cra_waitrequest
	wire   [63:0] acl_iface_kernel_cra_readdata;                                   // mm_interconnect_3:acl_iface_kernel_cra_readdata -> acl_iface:kernel_cra_readdata
	wire          acl_iface_kernel_cra_debugaccess;                                // acl_iface:kernel_cra_debugaccess -> mm_interconnect_3:acl_iface_kernel_cra_debugaccess
	wire   [29:0] acl_iface_kernel_cra_address;                                    // acl_iface:kernel_cra_address -> mm_interconnect_3:acl_iface_kernel_cra_address
	wire          acl_iface_kernel_cra_read;                                       // acl_iface:kernel_cra_read -> mm_interconnect_3:acl_iface_kernel_cra_read
	wire    [7:0] acl_iface_kernel_cra_byteenable;                                 // acl_iface:kernel_cra_byteenable -> mm_interconnect_3:acl_iface_kernel_cra_byteenable
	wire          acl_iface_kernel_cra_readdatavalid;                              // mm_interconnect_3:acl_iface_kernel_cra_readdatavalid -> acl_iface:kernel_cra_readdatavalid
	wire   [63:0] acl_iface_kernel_cra_writedata;                                  // acl_iface:kernel_cra_writedata -> mm_interconnect_3:acl_iface_kernel_cra_writedata
	wire          acl_iface_kernel_cra_write;                                      // acl_iface:kernel_cra_write -> mm_interconnect_3:acl_iface_kernel_cra_write
	wire    [0:0] acl_iface_kernel_cra_burstcount;                                 // acl_iface:kernel_cra_burstcount -> mm_interconnect_3:acl_iface_kernel_cra_burstcount
	wire   [63:0] mm_interconnect_3_cra_root_cra_slave_readdata;                   // cra_root:avs_readdata -> mm_interconnect_3:cra_root_cra_slave_readdata
	wire          mm_interconnect_3_cra_root_cra_slave_waitrequest;                // cra_root:avs_waitrequest -> mm_interconnect_3:cra_root_cra_slave_waitrequest
	wire    [3:0] mm_interconnect_3_cra_root_cra_slave_address;                    // mm_interconnect_3:cra_root_cra_slave_address -> cra_root:avs_addr
	wire          mm_interconnect_3_cra_root_cra_slave_read;                       // mm_interconnect_3:cra_root_cra_slave_read -> cra_root:avs_read
	wire    [7:0] mm_interconnect_3_cra_root_cra_slave_byteenable;                 // mm_interconnect_3:cra_root_cra_slave_byteenable -> cra_root:avs_byteena
	wire          mm_interconnect_3_cra_root_cra_slave_readdatavalid;              // cra_root:avs_readdatavalid -> mm_interconnect_3:cra_root_cra_slave_readdatavalid
	wire          mm_interconnect_3_cra_root_cra_slave_write;                      // mm_interconnect_3:cra_root_cra_slave_write -> cra_root:avs_write
	wire   [63:0] mm_interconnect_3_cra_root_cra_slave_writedata;                  // mm_interconnect_3:cra_root_cra_slave_writedata -> cra_root:avs_writedata
	wire          irq_mapper_receiver0_irq;                                        // genetic_algorithm_system:kernel_irq -> irq_mapper:receiver0_irq
	wire    [0:0] acl_iface_kernel_irq_irq;                                        // irq_mapper:sender_irq -> acl_iface:kernel_irq_irq
	wire          rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:acl_iface_global_reset_reset_bridge_in_reset_reset, mm_interconnect_0:acl_iface_kernel_mem0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:acl_iface_global_reset_reset_bridge_in_reset_reset, mm_interconnect_1:acl_iface_kernel_mem1_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_3:acl_iface_global_reset_reset_bridge_in_reset_reset, mm_interconnect_3:acl_iface_kernel_cra_translator_reset_reset_bridge_in_reset_reset]

	system_acl_iface acl_iface (
		.reset_n                               (global_reset_reset_n),                                  //               global_reset.reset_n
		.pcie_refclk_clk                       (pcie_refclk_clk),                                       //                pcie_refclk.clk
		.pcie_hip_serial_rx_in0                (pcie_rx_in0),                                           //            pcie_hip_serial.rx_in0
		.pcie_hip_serial_rx_in1                (pcie_rx_in1),                                           //                           .rx_in1
		.pcie_hip_serial_rx_in2                (pcie_rx_in2),                                           //                           .rx_in2
		.pcie_hip_serial_rx_in3                (pcie_rx_in3),                                           //                           .rx_in3
		.pcie_hip_serial_rx_in4                (pcie_rx_in4),                                           //                           .rx_in4
		.pcie_hip_serial_rx_in5                (pcie_rx_in5),                                           //                           .rx_in5
		.pcie_hip_serial_rx_in6                (pcie_rx_in6),                                           //                           .rx_in6
		.pcie_hip_serial_rx_in7                (pcie_rx_in7),                                           //                           .rx_in7
		.pcie_hip_serial_tx_out0               (pcie_tx_out0),                                          //                           .tx_out0
		.pcie_hip_serial_tx_out1               (pcie_tx_out1),                                          //                           .tx_out1
		.pcie_hip_serial_tx_out2               (pcie_tx_out2),                                          //                           .tx_out2
		.pcie_hip_serial_tx_out3               (pcie_tx_out3),                                          //                           .tx_out3
		.pcie_hip_serial_tx_out4               (pcie_tx_out4),                                          //                           .tx_out4
		.pcie_hip_serial_tx_out5               (pcie_tx_out5),                                          //                           .tx_out5
		.pcie_hip_serial_tx_out6               (pcie_tx_out6),                                          //                           .tx_out6
		.pcie_hip_serial_tx_out7               (pcie_tx_out7),                                          //                           .tx_out7
		.pcie_npor_npor                        (pcie_npor_npor),                                        //                  pcie_npor.npor
		.pcie_npor_pin_perst                   (pcie_npor_pin_perst),                                   //                           .pin_perst
		.ddr3a_mem_a                           (ddr3a_mem_a),                                           //                      ddr3a.mem_a
		.ddr3a_mem_ba                          (ddr3a_mem_ba),                                          //                           .mem_ba
		.ddr3a_mem_ck                          (ddr3a_mem_ck),                                          //                           .mem_ck
		.ddr3a_mem_ck_n                        (ddr3a_mem_ck_n),                                        //                           .mem_ck_n
		.ddr3a_mem_cke                         (ddr3a_mem_cke),                                         //                           .mem_cke
		.ddr3a_mem_cs_n                        (ddr3a_mem_cs_n),                                        //                           .mem_cs_n
		.ddr3a_mem_dm                          (ddr3a_mem_dm),                                          //                           .mem_dm
		.ddr3a_mem_ras_n                       (ddr3a_mem_ras_n),                                       //                           .mem_ras_n
		.ddr3a_mem_cas_n                       (ddr3a_mem_cas_n),                                       //                           .mem_cas_n
		.ddr3a_mem_we_n                        (ddr3a_mem_we_n),                                        //                           .mem_we_n
		.ddr3a_mem_reset_n                     (ddr3a_mem_reset_n),                                     //                           .mem_reset_n
		.ddr3a_mem_dq                          (ddr3a_mem_dq),                                          //                           .mem_dq
		.ddr3a_mem_dqs                         (ddr3a_mem_dqs),                                         //                           .mem_dqs
		.ddr3a_mem_dqs_n                       (ddr3a_mem_dqs_n),                                       //                           .mem_dqs_n
		.ddr3a_mem_odt                         (ddr3a_mem_odt),                                         //                           .mem_odt
		.octa_rzqin                            (ddr3a_mem_oct_rzqin),                                   //                       octa.rzqin
		.ddr3a_pll_ref_clk                     (ddr3a_pll_ref_clk),                                     //              ddr3a_pll_ref.clk
		.ddr3b_mem_a                           (ddr3b_mem_a),                                           //                      ddr3b.mem_a
		.ddr3b_mem_ba                          (ddr3b_mem_ba),                                          //                           .mem_ba
		.ddr3b_mem_ck                          (ddr3b_mem_ck),                                          //                           .mem_ck
		.ddr3b_mem_ck_n                        (ddr3b_mem_ck_n),                                        //                           .mem_ck_n
		.ddr3b_mem_cke                         (ddr3b_mem_cke),                                         //                           .mem_cke
		.ddr3b_mem_cs_n                        (ddr3b_mem_cs_n),                                        //                           .mem_cs_n
		.ddr3b_mem_dm                          (ddr3b_mem_dm),                                          //                           .mem_dm
		.ddr3b_mem_ras_n                       (ddr3b_mem_ras_n),                                       //                           .mem_ras_n
		.ddr3b_mem_cas_n                       (ddr3b_mem_cas_n),                                       //                           .mem_cas_n
		.ddr3b_mem_we_n                        (ddr3b_mem_we_n),                                        //                           .mem_we_n
		.ddr3b_mem_reset_n                     (ddr3b_mem_reset_n),                                     //                           .mem_reset_n
		.ddr3b_mem_dq                          (ddr3b_mem_dq),                                          //                           .mem_dq
		.ddr3b_mem_dqs                         (ddr3b_mem_dqs),                                         //                           .mem_dqs
		.ddr3b_mem_dqs_n                       (ddr3b_mem_dqs_n),                                       //                           .mem_dqs_n
		.ddr3b_mem_odt                         (ddr3b_mem_odt),                                         //                           .mem_odt
		.octb_rzqin                            (ddr3b_mem_oct_rzqin),                                   //                       octb.rzqin
		.ddr3b_pll_ref_clk                     (ddr3b_pll_ref_clk),                                     //              ddr3b_pll_ref.clk
		.pcie_hip_ctrl_test_in                 (),                                                      //              pcie_hip_ctrl.test_in
		.pcie_hip_ctrl_simu_mode_pipe          (),                                                      //                           .simu_mode_pipe
		.config_clk_clk                        (config_clk_clk),                                        //                 config_clk.clk
		.acl_internal_memorg_kernel_mode       (),                                                      // acl_internal_memorg_kernel.mode
		.kernel_clk2x_clk                      (acl_iface_kernel_clk2x_clk),                            //               kernel_clk2x.clk
		.kernel_pll_refclk_clk                 (kernel_pll_refclk_clk),                                 //          kernel_pll_refclk.clk
		.kernel_cra_waitrequest                (acl_iface_kernel_cra_waitrequest),                      //                 kernel_cra.waitrequest
		.kernel_cra_readdata                   (acl_iface_kernel_cra_readdata),                         //                           .readdata
		.kernel_cra_readdatavalid              (acl_iface_kernel_cra_readdatavalid),                    //                           .readdatavalid
		.kernel_cra_burstcount                 (acl_iface_kernel_cra_burstcount),                       //                           .burstcount
		.kernel_cra_writedata                  (acl_iface_kernel_cra_writedata),                        //                           .writedata
		.kernel_cra_address                    (acl_iface_kernel_cra_address),                          //                           .address
		.kernel_cra_write                      (acl_iface_kernel_cra_write),                            //                           .write
		.kernel_cra_read                       (acl_iface_kernel_cra_read),                             //                           .read
		.kernel_cra_byteenable                 (acl_iface_kernel_cra_byteenable),                       //                           .byteenable
		.kernel_cra_debugaccess                (acl_iface_kernel_cra_debugaccess),                      //                           .debugaccess
		.kernel_irq_irq                        (acl_iface_kernel_irq_irq),                              //                 kernel_irq.irq
		.kernel_mem0_waitrequest               (mm_interconnect_0_acl_iface_kernel_mem0_waitrequest),   //                kernel_mem0.waitrequest
		.kernel_mem0_readdata                  (mm_interconnect_0_acl_iface_kernel_mem0_readdata),      //                           .readdata
		.kernel_mem0_readdatavalid             (mm_interconnect_0_acl_iface_kernel_mem0_readdatavalid), //                           .readdatavalid
		.kernel_mem0_burstcount                (mm_interconnect_0_acl_iface_kernel_mem0_burstcount),    //                           .burstcount
		.kernel_mem0_writedata                 (mm_interconnect_0_acl_iface_kernel_mem0_writedata),     //                           .writedata
		.kernel_mem0_address                   (mm_interconnect_0_acl_iface_kernel_mem0_address),       //                           .address
		.kernel_mem0_write                     (mm_interconnect_0_acl_iface_kernel_mem0_write),         //                           .write
		.kernel_mem0_read                      (mm_interconnect_0_acl_iface_kernel_mem0_read),          //                           .read
		.kernel_mem0_byteenable                (mm_interconnect_0_acl_iface_kernel_mem0_byteenable),    //                           .byteenable
		.kernel_mem0_debugaccess               (mm_interconnect_0_acl_iface_kernel_mem0_debugaccess),   //                           .debugaccess
		.kernel_mem1_waitrequest               (mm_interconnect_1_acl_iface_kernel_mem1_waitrequest),   //                kernel_mem1.waitrequest
		.kernel_mem1_readdata                  (mm_interconnect_1_acl_iface_kernel_mem1_readdata),      //                           .readdata
		.kernel_mem1_readdatavalid             (mm_interconnect_1_acl_iface_kernel_mem1_readdatavalid), //                           .readdatavalid
		.kernel_mem1_burstcount                (mm_interconnect_1_acl_iface_kernel_mem1_burstcount),    //                           .burstcount
		.kernel_mem1_writedata                 (mm_interconnect_1_acl_iface_kernel_mem1_writedata),     //                           .writedata
		.kernel_mem1_address                   (mm_interconnect_1_acl_iface_kernel_mem1_address),       //                           .address
		.kernel_mem1_write                     (mm_interconnect_1_acl_iface_kernel_mem1_write),         //                           .write
		.kernel_mem1_read                      (mm_interconnect_1_acl_iface_kernel_mem1_read),          //                           .read
		.kernel_mem1_byteenable                (mm_interconnect_1_acl_iface_kernel_mem1_byteenable),    //                           .byteenable
		.kernel_mem1_debugaccess               (mm_interconnect_1_acl_iface_kernel_mem1_debugaccess),   //                           .debugaccess
		.acl_internal_snoop_data               (),                                                      //         acl_internal_snoop.data
		.acl_internal_snoop_valid              (),                                                      //                           .valid
		.acl_internal_snoop_ready              (),                                                      //                           .ready
		.kernel_clk_clk                        (acl_iface_kernel_clk_clk),                              //                 kernel_clk.clk
		.kernel_reset_reset_n                  (acl_iface_kernel_reset_reset),                          //               kernel_reset.reset_n
		.pcie_npor_out_reset_n                 (pcie_npor_out_reset_n),                                 //              pcie_npor_out.reset_n
		.reconfig_to_xcvr_reconfig_to_xcvr     (reconfig_to_xcvr_reconfig_to_xcvr),                     //           reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr_reconfig_from_xcvr (reconfig_from_xcvr_reconfig_from_xcvr)                  //         reconfig_from_xcvr.reconfig_from_xcvr
	);

	cra_ring_node #(
		.RING_ADDR_W (4),
		.CRA_ADDR_W  (4),
		.DATA_W      (64),
		.ID_W        (0),
		.ID          (32'b00000000000000000000000000000000)
	) avs_vadd_cra_cra_ring (
		.clk               (acl_iface_kernel_clk_clk),                       //      clock.clk
		.rst_n             (acl_iface_kernel_reset_reset),                   //      reset.reset_n
		.avm_read          (avs_vadd_cra_cra_ring_cra_master_read),          // cra_master.read
		.avm_write         (avs_vadd_cra_cra_ring_cra_master_write),         //           .write
		.avm_addr          (avs_vadd_cra_cra_ring_cra_master_address),       //           .address
		.avm_byteena       (avs_vadd_cra_cra_ring_cra_master_byteenable),    //           .byteenable
		.avm_writedata     (avs_vadd_cra_cra_ring_cra_master_writedata),     //           .writedata
		.avm_readdata      (avs_vadd_cra_cra_ring_cra_master_readdata),      //           .readdata
		.avm_readdatavalid (avs_vadd_cra_cra_ring_cra_master_readdatavalid), //           .readdatavalid
		.ri_read           (cra_root_ring_out_read),                         //    ring_in.read
		.ri_write          (cra_root_ring_out_write),                        //           .write
		.ri_addr           (cra_root_ring_out_addr),                         //           .addr
		.ri_data           (cra_root_ring_out_data),                         //           .data
		.ri_byteena        (cra_root_ring_out_byteena),                      //           .byteena
		.ri_datavalid      (cra_root_ring_out_datavalid),                    //           .datavalid
		.ro_read           (avs_vadd_cra_cra_ring_ring_out_read),            //   ring_out.read
		.ro_write          (avs_vadd_cra_cra_ring_ring_out_write),           //           .write
		.ro_addr           (avs_vadd_cra_cra_ring_ring_out_addr),            //           .addr
		.ro_data           (avs_vadd_cra_cra_ring_ring_out_data),            //           .data
		.ro_byteena        (avs_vadd_cra_cra_ring_ring_out_byteena),         //           .byteena
		.ro_datavalid      (avs_vadd_cra_cra_ring_ring_out_datavalid)        //           .datavalid
	);

	cra_ring_root #(
		.ADDR_W     (4),
		.DATA_W     (64),
		.ID_W       (0),
		.ROM_EXT_W  (0),
		.ROM_ENABLE (0)
	) cra_root (
		.clk               (acl_iface_kernel_clk_clk),                           //     clock.clk
		.rst_n             (acl_iface_kernel_reset_reset),                       //     reset.reset_n
		.avs_write         (mm_interconnect_3_cra_root_cra_slave_write),         // cra_slave.write
		.avs_addr          (mm_interconnect_3_cra_root_cra_slave_address),       //          .address
		.avs_byteena       (mm_interconnect_3_cra_root_cra_slave_byteenable),    //          .byteenable
		.avs_writedata     (mm_interconnect_3_cra_root_cra_slave_writedata),     //          .writedata
		.avs_readdata      (mm_interconnect_3_cra_root_cra_slave_readdata),      //          .readdata
		.avs_readdatavalid (mm_interconnect_3_cra_root_cra_slave_readdatavalid), //          .readdatavalid
		.avs_waitrequest   (mm_interconnect_3_cra_root_cra_slave_waitrequest),   //          .waitrequest
		.avs_read          (mm_interconnect_3_cra_root_cra_slave_read),          //          .read
		.ri_write          (avs_vadd_cra_cra_ring_ring_out_write),               //   ring_in.write
		.ri_addr           (avs_vadd_cra_cra_ring_ring_out_addr),                //          .addr
		.ri_byteena        (avs_vadd_cra_cra_ring_ring_out_byteena),             //          .byteena
		.ri_data           (avs_vadd_cra_cra_ring_ring_out_data),                //          .data
		.ri_read           (avs_vadd_cra_cra_ring_ring_out_read),                //          .read
		.ri_datavalid      (avs_vadd_cra_cra_ring_ring_out_datavalid),           //          .datavalid
		.ro_read           (cra_root_ring_out_read),                             //  ring_out.read
		.ro_write          (cra_root_ring_out_write),                            //          .write
		.ro_addr           (cra_root_ring_out_addr),                             //          .addr
		.ro_data           (cra_root_ring_out_data),                             //          .data
		.ro_byteena        (cra_root_ring_out_byteena),                          //          .byteena
		.ro_datavalid      (cra_root_ring_out_datavalid)                         //          .datavalid
	);

	genetic_algorithm_system genetic_algorithm_system (
		.clock                                  (acl_iface_kernel_clk_clk),                                        //              clock_reset.clk
		.resetn                                 (acl_iface_kernel_reset_reset),                                    //        clock_reset_reset.reset_n
		.clock2x                                (acl_iface_kernel_clk2x_clk),                                      //            clock_reset2x.clk
		.avs_vadd_cra_read                      (avs_vadd_cra_cra_ring_cra_master_read),                           //             avs_vadd_cra.read
		.avs_vadd_cra_write                     (avs_vadd_cra_cra_ring_cra_master_write),                          //                         .write
		.avs_vadd_cra_address                   (avs_vadd_cra_cra_ring_cra_master_address),                        //                         .address
		.avs_vadd_cra_writedata                 (avs_vadd_cra_cra_ring_cra_master_writedata),                      //                         .writedata
		.avs_vadd_cra_byteenable                (avs_vadd_cra_cra_ring_cra_master_byteenable),                     //                         .byteenable
		.avs_vadd_cra_readdata                  (avs_vadd_cra_cra_ring_cra_master_readdata),                       //                         .readdata
		.avs_vadd_cra_readdatavalid             (avs_vadd_cra_cra_ring_cra_master_readdatavalid),                  //                         .readdatavalid
		.kernel_irq                             (irq_mapper_receiver0_irq),                                        //               kernel_irq.irq
		.avm_memgmem0_port_0_0_rw_address       (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_address),       // avm_memgmem0_port_0_0_rw.address
		.avm_memgmem0_port_0_0_rw_read          (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_read),          //                         .read
		.avm_memgmem0_port_0_0_rw_write         (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_write),         //                         .write
		.avm_memgmem0_port_0_0_rw_writedata     (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_writedata),     //                         .writedata
		.avm_memgmem0_port_0_0_rw_byteenable    (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_byteenable),    //                         .byteenable
		.avm_memgmem0_port_0_0_rw_readdata      (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_readdata),      //                         .readdata
		.avm_memgmem0_port_0_0_rw_burstcount    (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_burstcount),    //                         .burstcount
		.avm_memgmem0_port_0_0_rw_waitrequest   (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_waitrequest),   //                         .waitrequest
		.avm_memgmem0_port_0_0_rw_readdatavalid (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_readdatavalid), //                         .readdatavalid
		.avm_memgmem0_port_1_0_rw_address       (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_address),       // avm_memgmem0_port_1_0_rw.address
		.avm_memgmem0_port_1_0_rw_read          (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_read),          //                         .read
		.avm_memgmem0_port_1_0_rw_write         (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_write),         //                         .write
		.avm_memgmem0_port_1_0_rw_writedata     (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_writedata),     //                         .writedata
		.avm_memgmem0_port_1_0_rw_byteenable    (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_byteenable),    //                         .byteenable
		.avm_memgmem0_port_1_0_rw_readdata      (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_readdata),      //                         .readdata
		.avm_memgmem0_port_1_0_rw_burstcount    (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_burstcount),    //                         .burstcount
		.avm_memgmem0_port_1_0_rw_waitrequest   (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_waitrequest),   //                         .waitrequest
		.avm_memgmem0_port_1_0_rw_readdatavalid (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_readdatavalid)  //                         .readdatavalid
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.acl_iface_kernel_clk_clk                                               (acl_iface_kernel_clk_clk),                                        //                                             acl_iface_kernel_clk.clk
		.acl_iface_global_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                                  //                     acl_iface_global_reset_reset_bridge_in_reset.reset
		.acl_iface_kernel_mem0_translator_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                                  //     acl_iface_kernel_mem0_translator_reset_reset_bridge_in_reset.reset
		.genetic_algorithm_system_clock_reset_reset_reset_bridge_in_reset_reset (~acl_iface_kernel_reset_reset),                                   // genetic_algorithm_system_clock_reset_reset_reset_bridge_in_reset.reset
		.genetic_algorithm_system_avm_memgmem0_port_0_0_rw_address              (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_address),       //                genetic_algorithm_system_avm_memgmem0_port_0_0_rw.address
		.genetic_algorithm_system_avm_memgmem0_port_0_0_rw_waitrequest          (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_waitrequest),   //                                                                 .waitrequest
		.genetic_algorithm_system_avm_memgmem0_port_0_0_rw_burstcount           (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_burstcount),    //                                                                 .burstcount
		.genetic_algorithm_system_avm_memgmem0_port_0_0_rw_byteenable           (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_byteenable),    //                                                                 .byteenable
		.genetic_algorithm_system_avm_memgmem0_port_0_0_rw_read                 (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_read),          //                                                                 .read
		.genetic_algorithm_system_avm_memgmem0_port_0_0_rw_readdata             (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_readdata),      //                                                                 .readdata
		.genetic_algorithm_system_avm_memgmem0_port_0_0_rw_readdatavalid        (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_readdatavalid), //                                                                 .readdatavalid
		.genetic_algorithm_system_avm_memgmem0_port_0_0_rw_write                (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_write),         //                                                                 .write
		.genetic_algorithm_system_avm_memgmem0_port_0_0_rw_writedata            (genetic_algorithm_system_avm_memgmem0_port_0_0_rw_writedata),     //                                                                 .writedata
		.acl_iface_kernel_mem0_address                                          (mm_interconnect_0_acl_iface_kernel_mem0_address),                 //                                            acl_iface_kernel_mem0.address
		.acl_iface_kernel_mem0_write                                            (mm_interconnect_0_acl_iface_kernel_mem0_write),                   //                                                                 .write
		.acl_iface_kernel_mem0_read                                             (mm_interconnect_0_acl_iface_kernel_mem0_read),                    //                                                                 .read
		.acl_iface_kernel_mem0_readdata                                         (mm_interconnect_0_acl_iface_kernel_mem0_readdata),                //                                                                 .readdata
		.acl_iface_kernel_mem0_writedata                                        (mm_interconnect_0_acl_iface_kernel_mem0_writedata),               //                                                                 .writedata
		.acl_iface_kernel_mem0_burstcount                                       (mm_interconnect_0_acl_iface_kernel_mem0_burstcount),              //                                                                 .burstcount
		.acl_iface_kernel_mem0_byteenable                                       (mm_interconnect_0_acl_iface_kernel_mem0_byteenable),              //                                                                 .byteenable
		.acl_iface_kernel_mem0_readdatavalid                                    (mm_interconnect_0_acl_iface_kernel_mem0_readdatavalid),           //                                                                 .readdatavalid
		.acl_iface_kernel_mem0_waitrequest                                      (mm_interconnect_0_acl_iface_kernel_mem0_waitrequest),             //                                                                 .waitrequest
		.acl_iface_kernel_mem0_debugaccess                                      (mm_interconnect_0_acl_iface_kernel_mem0_debugaccess)              //                                                                 .debugaccess
	);

	system_mm_interconnect_1 mm_interconnect_1 (
		.acl_iface_kernel_clk_clk                                               (acl_iface_kernel_clk_clk),                                        //                                             acl_iface_kernel_clk.clk
		.acl_iface_global_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                                  //                     acl_iface_global_reset_reset_bridge_in_reset.reset
		.acl_iface_kernel_mem1_translator_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                                  //     acl_iface_kernel_mem1_translator_reset_reset_bridge_in_reset.reset
		.genetic_algorithm_system_clock_reset_reset_reset_bridge_in_reset_reset (~acl_iface_kernel_reset_reset),                                   // genetic_algorithm_system_clock_reset_reset_reset_bridge_in_reset.reset
		.genetic_algorithm_system_avm_memgmem0_port_1_0_rw_address              (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_address),       //                genetic_algorithm_system_avm_memgmem0_port_1_0_rw.address
		.genetic_algorithm_system_avm_memgmem0_port_1_0_rw_waitrequest          (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_waitrequest),   //                                                                 .waitrequest
		.genetic_algorithm_system_avm_memgmem0_port_1_0_rw_burstcount           (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_burstcount),    //                                                                 .burstcount
		.genetic_algorithm_system_avm_memgmem0_port_1_0_rw_byteenable           (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_byteenable),    //                                                                 .byteenable
		.genetic_algorithm_system_avm_memgmem0_port_1_0_rw_read                 (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_read),          //                                                                 .read
		.genetic_algorithm_system_avm_memgmem0_port_1_0_rw_readdata             (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_readdata),      //                                                                 .readdata
		.genetic_algorithm_system_avm_memgmem0_port_1_0_rw_readdatavalid        (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_readdatavalid), //                                                                 .readdatavalid
		.genetic_algorithm_system_avm_memgmem0_port_1_0_rw_write                (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_write),         //                                                                 .write
		.genetic_algorithm_system_avm_memgmem0_port_1_0_rw_writedata            (genetic_algorithm_system_avm_memgmem0_port_1_0_rw_writedata),     //                                                                 .writedata
		.acl_iface_kernel_mem1_address                                          (mm_interconnect_1_acl_iface_kernel_mem1_address),                 //                                            acl_iface_kernel_mem1.address
		.acl_iface_kernel_mem1_write                                            (mm_interconnect_1_acl_iface_kernel_mem1_write),                   //                                                                 .write
		.acl_iface_kernel_mem1_read                                             (mm_interconnect_1_acl_iface_kernel_mem1_read),                    //                                                                 .read
		.acl_iface_kernel_mem1_readdata                                         (mm_interconnect_1_acl_iface_kernel_mem1_readdata),                //                                                                 .readdata
		.acl_iface_kernel_mem1_writedata                                        (mm_interconnect_1_acl_iface_kernel_mem1_writedata),               //                                                                 .writedata
		.acl_iface_kernel_mem1_burstcount                                       (mm_interconnect_1_acl_iface_kernel_mem1_burstcount),              //                                                                 .burstcount
		.acl_iface_kernel_mem1_byteenable                                       (mm_interconnect_1_acl_iface_kernel_mem1_byteenable),              //                                                                 .byteenable
		.acl_iface_kernel_mem1_readdatavalid                                    (mm_interconnect_1_acl_iface_kernel_mem1_readdatavalid),           //                                                                 .readdatavalid
		.acl_iface_kernel_mem1_waitrequest                                      (mm_interconnect_1_acl_iface_kernel_mem1_waitrequest),             //                                                                 .waitrequest
		.acl_iface_kernel_mem1_debugaccess                                      (mm_interconnect_1_acl_iface_kernel_mem1_debugaccess)              //                                                                 .debugaccess
	);

	system_mm_interconnect_3 mm_interconnect_3 (
		.acl_iface_kernel_clk_clk                                          (acl_iface_kernel_clk_clk),                           //                                        acl_iface_kernel_clk.clk
		.acl_iface_global_reset_reset_bridge_in_reset_reset                (rst_controller_reset_out_reset),                     //                acl_iface_global_reset_reset_bridge_in_reset.reset
		.acl_iface_kernel_cra_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                     // acl_iface_kernel_cra_translator_reset_reset_bridge_in_reset.reset
		.cra_root_reset_reset_bridge_in_reset_reset                        (~acl_iface_kernel_reset_reset),                      //                        cra_root_reset_reset_bridge_in_reset.reset
		.acl_iface_kernel_cra_address                                      (acl_iface_kernel_cra_address),                       //                                        acl_iface_kernel_cra.address
		.acl_iface_kernel_cra_waitrequest                                  (acl_iface_kernel_cra_waitrequest),                   //                                                            .waitrequest
		.acl_iface_kernel_cra_burstcount                                   (acl_iface_kernel_cra_burstcount),                    //                                                            .burstcount
		.acl_iface_kernel_cra_byteenable                                   (acl_iface_kernel_cra_byteenable),                    //                                                            .byteenable
		.acl_iface_kernel_cra_read                                         (acl_iface_kernel_cra_read),                          //                                                            .read
		.acl_iface_kernel_cra_readdata                                     (acl_iface_kernel_cra_readdata),                      //                                                            .readdata
		.acl_iface_kernel_cra_readdatavalid                                (acl_iface_kernel_cra_readdatavalid),                 //                                                            .readdatavalid
		.acl_iface_kernel_cra_write                                        (acl_iface_kernel_cra_write),                         //                                                            .write
		.acl_iface_kernel_cra_writedata                                    (acl_iface_kernel_cra_writedata),                     //                                                            .writedata
		.acl_iface_kernel_cra_debugaccess                                  (acl_iface_kernel_cra_debugaccess),                   //                                                            .debugaccess
		.cra_root_cra_slave_address                                        (mm_interconnect_3_cra_root_cra_slave_address),       //                                          cra_root_cra_slave.address
		.cra_root_cra_slave_write                                          (mm_interconnect_3_cra_root_cra_slave_write),         //                                                            .write
		.cra_root_cra_slave_read                                           (mm_interconnect_3_cra_root_cra_slave_read),          //                                                            .read
		.cra_root_cra_slave_readdata                                       (mm_interconnect_3_cra_root_cra_slave_readdata),      //                                                            .readdata
		.cra_root_cra_slave_writedata                                      (mm_interconnect_3_cra_root_cra_slave_writedata),     //                                                            .writedata
		.cra_root_cra_slave_byteenable                                     (mm_interconnect_3_cra_root_cra_slave_byteenable),    //                                                            .byteenable
		.cra_root_cra_slave_readdatavalid                                  (mm_interconnect_3_cra_root_cra_slave_readdatavalid), //                                                            .readdatavalid
		.cra_root_cra_slave_waitrequest                                    (mm_interconnect_3_cra_root_cra_slave_waitrequest)    //                                                            .waitrequest
	);

	system_irq_mapper irq_mapper (
		.clk           (acl_iface_kernel_clk_clk),       //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (acl_iface_kernel_irq_irq)        //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~global_reset_reset_n),          // reset_in0.reset
		.clk            (acl_iface_kernel_clk_clk),       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
